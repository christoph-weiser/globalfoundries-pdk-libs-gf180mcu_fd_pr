* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

*******************************************************************************
* Document No.      : YI-141-SM064
* Revision          : 9
* Process Name      : 0.18um 3.3V/6V high voltage MCU process
* Process ID        : TH18300G0A-PID007347
*					  TH18300G1A-PID007352
*					  TH183G0G6A-PID009507
*					  TH18300G7A-PID009628
*					  TH18300G4A-PID009792
*					  TH18300G9A-PID010186
* Wafer ID          : GT3512K wf#02 (3.3V NMOS, 6.0V NMOS, 6.0V native NMOS and NMOSCAP)
*                     GT3512K wf#06 (3.3V PMOS, 6.0V PMOS, PMOSCAP and BJT)
*                     GT9755L wf#18 (PWELL/DNWELL and DNWELL/Psub diode, Vertical NPN)
*                     JT1042L01 (6V NMOS L=0.6um)
*                     TCXN39W20 W#4 schottky diode
************************************************************************************************
* Models included in this release :
*
*      ModelName          Description
*      ---------          -----------
*      nmos_3p3           Subcircuit model for 3.3V NMOS
*      pmos_3p3           Subcircuit model for 3.3V PMOS
*      nmos_6p0           Subcircuit model for 6.0V NMOS
*      pmos_6p0           Subcircuit model for 6.0V PMOS
*      nmos_3p3_sab       Subcircuit model for 3.3V NMOS with Drain side SAB
*      pmos_3p3_sab       Subcircuit model for 3.3V PMOS with Drain side SAB
*      nmos_6p0_sab       Subcircuit model for 6.0V NMOS with Drain side SAB
*      pmos_6p0_sab       Subcircuit model for 6.0V PMOS with Drain side SAB
*      nmos_6p0_nat       Subcircuit model for 6.0V native NMOS
*
*      np_3p3             Model for 3.3V N+/Psub diode
*      pn_3p3             Model for 3.3V P+/Nwell diode
*      np_6p0             Model for 6.0V N+/Psub diode
*      pn_6p0             Model for 6.0V P+/Nwell diode
*      nwp_3p3            Model for 3.3V Nwell/Psub diode
*      nwp_6p0            Model for 6.0V Nwell/Psub diode
*      dnwpw              Model for PWELL/DNWELL diode
*      dnwps	          Model for DNWELL/Psub diode
*      sc_diode           Model for Schottky Diode
*
*      vpnp_0p42x10       Subcircuit GP model for VPNP with emitter size of 10umx0.42um
*      vpnp_0p42x5        Subcircuit GP model for VPNP with emitter size of 5umx0.42um
*      vpnp_10x10         Subcircuit GP model for VPNP with emitter size of 10umx10um
*      vpnp_5x5           Subcircuit GP model for VPNP with emitter size of 5umx5um
*      vnpn_10x10         Subcircuit GP model for VNPN with emitter size of 10umx10um(four terminal)
*      vnpn_5x5        	  Subcircuit GP model for VNPN with emitter size of 5umx5um(four terminal)
*      vnpn_0p54x16       Subcircuit GP model for VNPN with emitter size of 0.54umx16um(four terminal)
*      vnpn_0p54x8        Subcircuit GP model for VNPN with emitter size of 0.54umx8um(four terminal)
*      vnpn_0p54x4        Subcircuit GP model for VNPN with emitter size of 0.54umx4um(four terminal)
*      vnpn_0p54x2        Subcircuit GP model for VNPN with emitter size of 0.54umx2um(four terminal)
*
*      nplus_u            Subcircuit Model for 3-terminal unsalicided n+ diffusion resistor
*      pplus_u            Subcircuit Model for 3-terminal unsalicided P+ diffusion resistor
*      nplus_s            Subcircuit Model for 3-terminal salicided N+ diffusion resistor
*      pplus_s            Subcircuit Model for 3-terminal salicided P+ diffusion resistor
*      nwell              Subcircuit Model for 3-terminal nwell resistor under STI
*      npolyf_u           Subcircuit Model for 3-terminal unsalicided n+ poly resistor
*      ppolyf_u           Subcircuit Model for 3-terminal unsalicided p+ poly resistor
*      npolyf_s           Subcircuit Model for 3-terminal salicided n+ poly resistor
*      ppolyf_s           Subcircuit Model for 3-terminal salicided p+ poly resistor
*      ppolyf_u_1k        Subcircuit Model for 3-terminal 1k high-Rs p+ poly resistor on field oxide (3.3V area)
*      ppolyf_u_2k        Subcircuit Model for 3-terminal 2k high-Rs p+ poly resistor on field oxide (3.3V area)
*      ppolyf_u_1k_6p0    Subcircuit Model for 3-terminal 1k high-Rs p+ poly resistor on field oxide (6.0V area)
*      ppolyf_u_2k_6p0    Subcircuit Model for 3-terminal 2k high-Rs p+ poly resistor on field oxide (6.0V area)
*      ppolyf_u_3k        Subcircuit Model for 3-terminal 3k high-Rs p+ poly resistor on field oxide (both 3.3V & 6.0V area)
*      rm1                Subcircuit Model for 2-terminal metal 1 resistor
*      rm2                Subcircuit Model for 2-terminal metal 2 resistor
*      rm3                Subcircuit Model for 2-terminal metal 3 resistor
*      tm6k               Subcircuit Model for 2-terminal top metal 6k resistor
*      tm9k               Subcircuit Model for 2-terminal top metal 9k resistor
*      tm11k              Subcircuit Model for 2-terminal top metal 11k resistor
*      tm30k              Subcircuit Model for 2-terminal top metal 30k resistor
*
*      mim_1p5fF          Subcircuit Model for 1.5fF/um2 MIM (*)-usable for Volt <=6V across capacitor
*      mim_1p0fF          Subcircuit Model for 1.0fF/um2 MIM (*)-usable for Volt <=20V across capacitor
*      mim_2p0fF          Subcircuit Model for 2fF/um2 MIM      -usable for Volt <=6V across capacitor
*
*      nmoscap_3p3        Subcircuit Model for 3.3v inversion-mode  NMOS capacitor
*      pmoscap_3p3	 	  Subcircuit Model for 3.3v inversion-mode  PMOS capacitor
*      nmoscap_6p0        Subcircuit Model for 6.0V inversion-mode  NMOS capacitor
*      pmoscap_6p0	  	  Subcircuit Model for 6.0V inversion-mode  PMOS capacitor
*      nmoscap_3p3_b      Subcircuit Model for 3.3v NMOS in Nwell capacitor
*      pmoscap_3p3_b	  Subcircuit Model for 3.3v PMOS in Pwell capacitor
*      nmoscap_6p0_b      Subcircuit Model for 6.0V NMOS in Nwell capacitor
*      pmoscap_6p0_b	  Subcircuit Model for 6.0V PMOS in Pwell capacitor
*
*      efuse    	      Subcircuit model for 6V/(5V) efuse
************************************************************************************************

.options parser model_binning=true

.lib typical
.lib 'sm141064.spice' nmos_3p3_t
.lib 'sm141064.spice' pmos_3p3_t
.param rsh_nplus_u_m=60
.param rsh_pplus_u_m=185
.param nmos_6p0_vsat=1
.param nmos_6p0_vth0=0
.param nmos_6p0_xl=0
.param nmos_6p0_xw=0
.param nmos_6p0_tox=0
.param nmos_6p0_cgso=1
.param nmos_6p0_cgdo=1
.param nmos_6p0_nat_u0='0.070102'
.param nmos_6p0_nat_vth0='-0.039'
.param nmos_6p0_nat_xl='0'
.param nmos_6p0_nat_xw='0'
.param nmos_6p0_nat_tox='1.52e-008'
.param nmos_6p0_nat_cgso='1e-010'
.param nmos_6p0_nat_cgdo='1e-010'
.param pmos_6p0_dvth0=0
.param pmos_6p0_dxl=0
.param pmos_6p0_dxw=0
.param pmos_6p0_dtox=0
.param pmos_6p0_dcgdo=1
.param pmos_6p0_dcgso=1
.lib 'sm141064.spice' nmos_6p0_t
.lib 'sm141064.spice' pmos_6p0_t
.lib 'sm141064.spice' nmos_6p0_nat_t
.lib 'sm141064.spice' noise_corner
.lib 'sm141064.spice' fets_mm
.endl typical

.lib ff
.lib 'sm141064.spice' nmos_3p3_f
.lib 'sm141064.spice' pmos_3p3_f
.param rsh_nplus_u_m=45
.param rsh_pplus_u_m=145
.param nmos_6p0_vsat=1.0846
.param nmos_6p0_vth0=-0.1298
.param nmos_6p0_xl=-4.2e-8
.param nmos_6p0_xw=5e-8
.param nmos_6p0_tox=-1e-9
.param nmos_6p0_cgso=0.9
.param nmos_6p0_cgdo=0.9
.param nmos_6p0_nat_u0='0.118'
.param nmos_6p0_nat_vth0='-0.216'
.param nmos_6p0_nat_xl='-2e-7'
.param nmos_6p0_nat_xw='1e-7'
.param nmos_6p0_nat_tox='1.42e-008'
.param nmos_6p0_nat_cgso='9e-011'
.param nmos_6p0_nat_cgdo='9e-011'
.param pmos_6p0_dvth0=0.1245
.param pmos_6p0_dxl=-4.65e-8
.param pmos_6p0_dxw=5e-8
.param pmos_6p0_dtox=-1e-9
.param pmos_6p0_dcgdo=0.9
.param pmos_6p0_dcgso=0.9
.lib 'sm141064.spice' nmos_6p0_t
.lib 'sm141064.spice' pmos_6p0_t
.lib 'sm141064.spice' nmos_6p0_nat_t
.lib 'sm141064.spice' noise_corner
.lib 'sm141064.spice' fets_mm
.endl ff

.lib ss
.lib 'sm141064.spice' nmos_3p3_s
.lib 'sm141064.spice' pmos_3p3_s
.param rsh_nplus_u_m=75
.param rsh_pplus_u_m=225
.param nmos_6p0_vsat=0.899
.param nmos_6p0_vth0=0.1193
.param nmos_6p0_xl=7e-8
.param nmos_6p0_xw=-5e-8
.param nmos_6p0_tox=1e-9
.param nmos_6p0_cgso=1.1
.param nmos_6p0_cgdo=1.1
.param nmos_6p0_nat_u0='0.046'
.param nmos_6p0_nat_vth0='0.1417'
.param nmos_6p0_nat_xl='2e-7'
.param nmos_6p0_nat_xw='-1e-7'
.param nmos_6p0_nat_tox='1.62e-008'
.param nmos_6p0_nat_cgso='1.1e-010'
.param nmos_6p0_nat_cgdo='1.1e-010'
.param pmos_6p0_dvth0=-0.1225
.param pmos_6p0_dxl=6.9e-8
.param pmos_6p0_dxw=-5e-8
.param pmos_6p0_dtox=1e-9
.param pmos_6p0_dcgdo=1.1
.param pmos_6p0_dcgso=1.1
.lib 'sm141064.spice' nmos_6p0_t
.lib 'sm141064.spice' pmos_6p0_t
.lib 'sm141064.spice' nmos_6p0_nat_t
.lib 'sm141064.spice' noise_corner
.lib 'sm141064.spice' fets_mm
.endl ss

.lib fs
.lib 'sm141064.spice' nmos_3p3_fs
.lib 'sm141064.spice' pmos_3p3_fs
.param rsh_nplus_u_m=48
.param rsh_pplus_u_m=219
.param nmos_6p0_vsat='0.0846*0.67+1'
.param nmos_6p0_vth0='-0.1298*0.75'
.param nmos_6p0_xl='-4.2e-8*0.67'
.param nmos_6p0_xw='5e-8*0.67'
.param nmos_6p0_tox='-1e-9*0.75'
.param nmos_6p0_cgso=0.93
.param nmos_6p0_cgdo=0.93
.param nmos_6p0_nat_u0='0.102034'
.param nmos_6p0_nat_vth0='-0.157'
.param nmos_6p0_nat_xl='-1.33e-7'
.param nmos_6p0_nat_xw='6.7e-8'
.param nmos_6p0_nat_tox='1.453e-008'
.param nmos_6p0_nat_cgso='9.33e-011'
.param nmos_6p0_nat_cgdo='9.33e-011'
.param pmos_6p0_dvth0=-0.0829
.param pmos_6p0_dxl=4.1e-8
.param pmos_6p0_dxw=-3.35e-8
.param pmos_6p0_dtox=6.7e-10
.param pmos_6p0_dcgdo=1.07
.param pmos_6p0_dcgso=1.07
.lib 'sm141064.spice' nmos_6p0_t
.lib 'sm141064.spice' pmos_6p0_t
.lib 'sm141064.spice' nmos_6p0_nat_t
.lib 'sm141064.spice' noise_corner
.lib 'sm141064.spice' fets_mm
.endl fs

.lib sf
.lib 'sm141064.spice' nmos_3p3_sf
.lib 'sm141064.spice' pmos_3p3_sf
.param rsh_nplus_u_m=72
.param rsh_pplus_u_m=150
.param nmos_6p0_vsat='1-(1-0.899)*0.67'
.param nmos_6p0_vth0='0.1193*0.75'
.param nmos_6p0_xl='7e-8*0.67'
.param nmos_6p0_xw='-5e-8*0.67'
.param nmos_6p0_tox='1e-9*0.75'
.param nmos_6p0_cgso=1.07
.param nmos_6p0_cgdo=1.07
.param nmos_6p0_nat_u0='0.054034'
.param nmos_6p0_nat_vth0='0.08147'
.param nmos_6p0_nat_xl='1.33e-7'
.param nmos_6p0_nat_xw='-6.7e-8'
.param nmos_6p0_nat_tox='1.587e-008'
.param nmos_6p0_nat_cgso='1.067e-010'
.param nmos_6p0_nat_cgdo='1.067e-010'
.param pmos_6p0_dvth0=0.0827
.param pmos_6p0_dxl=-3.22e-8
.param pmos_6p0_dxw=3.35e-8
.param pmos_6p0_dtox=-6.7e-10
.param pmos_6p0_dcgdo=0.93
.param pmos_6p0_dcgso=0.93
.lib 'sm141064.spice' nmos_6p0_t
.lib 'sm141064.spice' pmos_6p0_t
.lib 'sm141064.spice' nmos_6p0_nat_t
.lib 'sm141064.spice' noise_corner
.lib 'sm141064.spice' fets_mm
.endl sf

.lib bjt_typical
.param isa=1
.param bfa=1
.param rba=1
.param rea=1
.param rca=1
.param rbma=1
.param cjea=1
.param cjca=1
.param is_cor_npn=1
.param bf_cor_npn=1
.param rb_cor_npn=1
.param re_cor_npn=1
.param rc_cor_npn=1
.param rbm_cor_npn=1
.param cjc_cor_npn=1
.param cje_cor_npn=1
.param mc_xis_vnpn=0
.param mc_xbf_vnpn=0
.param mc_xrb_vnpn=0
.param mc_xre_vnpn=0
.param mc_xrc_vnpn=0
.param mc_xcje_vnpn=0
.param mc_xcjc_vnpn=0
.param mc_xis_vpnp=0
.param mc_xbf_vpnp=0
.param mc_xrb_vpnp=0
.param mc_xre_vpnp=0
.param mc_xrc_vpnp=0
.param mc_xcje_vpnp=0
.param mc_xcjc_vpnp=0
.lib 'sm141064.spice' bjt_mc
.endl bjt_typical

.lib bjt_ss
.param isa=0.65
.param bfa=0.80
.param rba=1.2
.param rea=1.2
.param rca=1.2
.param rbma=1.2
.param cjea=1.15
.param cjca=1.15
.param is_cor_npn=0.4
.param bf_cor_npn=0.57
.param rb_cor_npn=1.2
.param re_cor_npn=1.2
.param rc_cor_npn=1.2
.param rbm_cor_npn=1.2
.param cjc_cor_npn=1.15
.param cje_cor_npn=1.15
.param mc_xis_vnpn=0
.param mc_xbf_vnpn=0
.param mc_xrb_vnpn=0
.param mc_xre_vnpn=0
.param mc_xrc_vnpn=0
.param mc_xcje_vnpn=0
.param mc_xcjc_vnpn=0
.param mc_xis_vpnp=0
.param mc_xbf_vpnp=0
.param mc_xrb_vpnp=0
.param mc_xre_vpnp=0
.param mc_xrc_vpnp=0
.param mc_xcje_vpnp=0
.param mc_xcjc_vpnp=0
.lib 'sm141064.spice' bjt_mc
.endl bjt_ss

.lib bjt_ff
.param isa=1.35
.param bfa=1.2
.param rba=0.8
.param rea=0.8
.param rca=0.8
.param rbma=0.8
.param cjea=0.85
.param cjca=0.85
.param is_cor_npn=2.25
.param bf_cor_npn=1.31
.param rb_cor_npn=0.8
.param re_cor_npn=0.8
.param rc_cor_npn=0.8
.param rbm_cor_npn=0.8
.param cjc_cor_npn=0.85
.param cje_cor_npn=0.85
.param mc_xis_vnpn=0
.param mc_xbf_vnpn=0
.param mc_xrb_vnpn=0
.param mc_xre_vnpn=0
.param mc_xrc_vnpn=0
.param mc_xcje_vnpn=0
.param mc_xcjc_vnpn=0
.param mc_xis_vpnp=0
.param mc_xbf_vpnp=0
.param mc_xrb_vpnp=0
.param mc_xre_vpnp=0
.param mc_xrc_vpnp=0
.param mc_xcje_vpnp=0
.param mc_xcjc_vpnp=0
.lib 'sm141064.spice' bjt_mc
.endl bjt_ff

.lib diode_typical
.param jsa=1
.param rsa=1
.param cja=1
.param cjswa=1
.param jsa_sc=0
.param vba_sc=0
.param rs_sc=1
.param jtuna_sc=0
.param cja_sc=1
.lib 'sm141064.spice' dio
.endl diode_typical

.lib diode_ss
.param jsa=0.85
.param rsa=1.1
.param cja=1.1
.param cjswa=1.1
.param jsa_sc=-1.6
.param vba_sc=-7
.param rs_sc=1.1
.param jtuna_sc=-0.77
.param cja_sc=1.1
.lib 'sm141064.spice' dio
.endl diode_ss

.lib diode_ff
.param jsa=1.15
.param rsa=0.9
.param cja=0.9
.param cjswa=0.9
.param jsa_sc=1.6
.param vba_sc=7
.param rs_sc=0.9
.param jtuna_sc=0.77
.param cja_sc=0.9
.lib 'sm141064.spice' dio
.endl diode_ff

.lib res_typical
.param rsh_nplus_u=60
.param rsh_pplus_u=185
.param rsh_nplus_s=6.3
.param rsh_pplus_s=7
.param rsh_nwell=1000
.param rsh_npolyf_u=310
.param rsh_ppolyf_u=350
.param rsh_npolyf_s=6.8
.param rsh_ppolyf_s=7.3
.param rsh_ppolyf_u_1k=1000
.param rsh_ppolyf_u_2k=2000
.param rsh_ppolyf_u_1k_6p0=1000
.param rsh_ppolyf_u_2k_6p0=2000
.param rsh_ppolyf_u_3k=3000
.param rsh_rm1=0.09
.param rsh_rm2=0.09
.param rsh_rm3=0.09
.param rsh_tm6k=60e-3
.param rsh_tm9k=40e-3
.param rsh_tm11k=40e-3
.param rsh_tm30k=9.5e-3
.lib 'sm141064.spice' res
.lib 'sm141064.spice' efuse
.lib 'sm141064.spice' res_statistical_par
.endl res_typical

.lib res_ss
.param rsh_nplus_u=75
.param rsh_pplus_u=225
.param rsh_nplus_s=15
.param rsh_pplus_s=15
.param rsh_nwell=1200
.param rsh_npolyf_u=370
.param rsh_ppolyf_u=420
.param rsh_npolyf_s=15
.param rsh_ppolyf_s=15
.param rsh_ppolyf_u_1k='1000+200'
.param rsh_ppolyf_u_2k='2000+400'
.param rsh_ppolyf_u_1k_6p0='1000+200'
.param rsh_ppolyf_u_2k_6p0='2000+400'
.param rsh_ppolyf_u_3k='3000+750'
.param rsh_rm1='0.09+0.012'
.param rsh_rm2='0.09+0.012'
.param rsh_rm3='0.09+0.012'
.param rsh_tm6k='60e-3+10e-3'
.param rsh_tm9k='40e-3+9e-3'
.param rsh_tm11k='40e-3+9e-3'
.param rsh_tm30k='9.5e-3+4.5e-3'
.lib 'sm141064.spice' res
.lib 'sm141064.spice' efuse
.lib 'sm141064.spice' res_statistical_par
.endl res_ss

.lib res_ff
.param rsh_nplus_u=45
.param rsh_pplus_u=145
.param rsh_nplus_s=1
.param rsh_pplus_s=1
.param rsh_nwell=800
.param rsh_npolyf_u=250
.param rsh_ppolyf_u=280
.param rsh_npolyf_s=1
.param rsh_ppolyf_s=1
.param rsh_ppolyf_u_1k='1000-200'
.param rsh_ppolyf_u_2k='2000-400'
.param rsh_ppolyf_u_1k_6p0='1000-200'
.param rsh_ppolyf_u_2k_6p0='2000-400'
.param rsh_ppolyf_u_3k='3000-750'
.param rsh_rm1='0.09-0.012'
.param rsh_rm2='0.09-0.012'
.param rsh_rm3='0.09-0.012'
.param rsh_tm6k='60e-3-10e-3'
.param rsh_tm9k='40e-3-9e-3'
.param rsh_tm11k='40e-3-9e-3'
.param rsh_tm30k='9.5e-3-3.5e-3'
.lib 'sm141064.spice' res
.lib 'sm141064.spice' efuse
.lib 'sm141064.spice' res_statistical_par
.endl res_ff

.lib mimcap_typical
.param mim_corner_1p5ff=1
.param mim_corner_1p0ff=1
.param mim_corner_2p0ff=1
.param mc_c_cox_1p0ff=0
.param mc_c_cox_1p5ff=0
.param mc_c_cox_2p0ff=0
.lib 'sm141064.spice' mim_cap
.endl mimcap_typical

.lib mimcap_ss
.param mim_corner_1p5ff=1.155
.param mim_corner_1p0ff=1.1
.param mim_corner_2p0ff=1.1
.param mc_c_cox_1p0ff=0
.param mc_c_cox_1p5ff=0
.param mc_c_cox_2p0ff=0
.lib 'sm141064.spice' mim_cap
.endl mimcap_ss

.lib mimcap_ff
.param mim_corner_1p5ff=0.845
.param mim_corner_1p0ff=0.9
.param mim_corner_2p0ff=0.9
.param mc_c_cox_1p0ff=0
.param mc_c_cox_1p5ff=0
.param mc_c_cox_2p0ff=0
.lib 'sm141064.spice' mim_cap
.endl mimcap_ff

.lib moscap_typical
.param nmoscap_3p3_corner=1
.param pmoscap_3p3_corner=1
.param nmoscap_6p0_corner=1
.param pmoscap_6p0_corner=1
.param nmoscap_3p3_b_corner=1
.param pmoscap_3p3_b_corner=1
.param nmoscap_6p0_b_corner=1
.param pmoscap_6p0_b_corner=1
.lib 'sm141064.spice' moscap
.endl moscap_typical

.lib moscap_ff
.param nmoscap_3p3_corner=0.9
.param pmoscap_3p3_corner=0.9
.param nmoscap_6p0_corner=0.9
.param pmoscap_6p0_corner=0.9
.param nmoscap_3p3_b_corner=0.9
.param pmoscap_3p3_b_corner=0.9
.param nmoscap_6p0_b_corner=0.9
.param pmoscap_6p0_b_corner=0.9
.lib 'sm141064.spice' moscap
.endl moscap_ff

.lib moscap_ss
.param nmoscap_3p3_corner=1.1
.param pmoscap_3p3_corner=1.1
.param nmoscap_6p0_corner=1.1
.param pmoscap_6p0_corner=1.1
.param nmoscap_3p3_b_corner=1.1
.param pmoscap_3p3_b_corner=1.1
.param nmoscap_6p0_b_corner=1.1
.param pmoscap_6p0_b_corner=1.1
.lib 'sm141064.spice' moscap
.endl moscap_ss

.lib statistical
.param mc_sig_vth2='agauss(0,1,3)'
.param mc_toxe2='agauss(0,1,3)'
.param mc_xl2='agauss(0,1,3)'
.param mc_xw2='agauss(0,1,3)'
.param mc_xj2='agauss(0,1,3)'
.param mc_sig_vthn2='agauss(0,1,3)'
.param mc_toxen2='agauss(0,1,3)'
.param mc_xln2='agauss(0,1,3)'
.param mc_xwn2='agauss(0,1,3)'
.param mc_xjn2='agauss(0,1,3)'
.param mc_rdswn2='agauss(0,1,3)'
.param mc_sig_vthp2='agauss(0,1,3)'
.param mc_toxep2='agauss(0,1,3)'
.param mc_xlp2='agauss(0,1,3)'
.param mc_xwp2='agauss(0,1,3)'
.param mc_xjp2='agauss(0,1,3)'
.param mc_rdswp2='agauss(0,1,3)'
.param mc_rsh_nplus_u_temp='agauss(0,3.85,3)'
.param mc_rsh_pplus_u_temp='agauss(0,10,3)'
.param mc_sig_vth='mc_sig_vth2'
.param mc_toxe='mc_toxe2'
.param mc_xl='mc_xl2'
.param mc_xw='mc_xw2'
.param mc_xj='mc_xj2'
.param mc_sig_vthn='mc_sig_vthn2'
.param mc_toxen='mc_toxen2'
.param mc_xln='mc_xln2'
.param mc_xwn='mc_xwn2'
.param mc_xjn='mc_xjn2'
.param mc_rdswn='mc_rdswn2'
.param mc_sig_vthp='mc_sig_vthp2'
.param mc_toxep='mc_toxep2'
.param mc_xlp='mc_xlp2'
.param mc_xwp='mc_xwp2'
.param mc_xjp='mc_xjp2'
.param mc_rdswp='mc_rdswp2'
.param mc_rsh_nplus_u='mc_rsh_nplus_u_temp'
.param mc_rsh_pplus_u='mc_rsh_pplus_u_temp'
.param nmos_3p3_sig_vth1='(5e-3*mc_sig_vth+30e-3*mc_sig_vthn)*sw_stat_global*mc_skew'
.param nmos_3p3_sig_vth2='(5e-3*mc_sig_vth+25e-3*mc_sig_vthn)*sw_stat_global*mc_skew'
.param nmos_3p3_sig_vth3='(5e-3*mc_sig_vth+15e-3*mc_sig_vthn)*sw_stat_global*mc_skew'
.param nmos_3p3_tox='8e-009+(1.6e-10*mc_toxe+0.3e-10*mc_toxen)*sw_stat_global*mc_skew'
.param nmos_3p3_xl='(7e-9*mc_xl+6e-9*mc_xln)*sw_stat_global*mc_skew'
.param nmos_3p3_xw='(7e-9*mc_xw+3e-9*mc_xwn)*sw_stat_global*mc_skew'
.param nmos_3p3_xj='1e-7+(0.3e-9*mc_xj+0.7e-9*mc_xjn)*sw_stat_global*mc_skew'
.param nmos_3p3_rdsw='530*(1+0.15*mc_rdswn*sw_stat_global*mc_skew)'
.param nmos_3p3_vth0_0='0.70837662+nmos_3p3_sig_vth1'
.param nmos_3p3_vth0_1='0.67781184+nmos_3p3_sig_vth1'
.param nmos_3p3_vth0_2='0.66097097+nmos_3p3_sig_vth2'
.param nmos_3p3_vth0_3='0.66064857+nmos_3p3_sig_vth2'
.param nmos_3p3_vth0_4='0.72356597+nmos_3p3_sig_vth1'
.param nmos_3p3_vth0_5='0.67504024+nmos_3p3_sig_vth2'
.param nmos_3p3_vth0_6='0.64923469+nmos_3p3_sig_vth2'
.param nmos_3p3_vth0_7='0.65055971+nmos_3p3_sig_vth3'
.param nmos_3p3_vth0_8='0.75419347+nmos_3p3_sig_vth2'
.param nmos_3p3_vth0_9='0.66260505+nmos_3p3_sig_vth2'
.param nmos_3p3_vth0_10='0.64815901+nmos_3p3_sig_vth3'
.param nmos_3p3_vth0_11='0.64889718+nmos_3p3_sig_vth3'
.param nmos_3p3_vth0_12='0.74840818+nmos_3p3_sig_vth2'
.param nmos_3p3_vth0_13='0.66297571+nmos_3p3_sig_vth3'
.param nmos_3p3_vth0_14='0.64787864+nmos_3p3_sig_vth3'
.param nmos_3p3_vth0_15='0.64857+nmos_3p3_sig_vth3'
.param pmos_3p3_sig_vth1='(-5e-3*mc_sig_vth-38e-3*mc_sig_vthp)*sw_stat_global*mc_skew'
.param pmos_3p3_sig_vth2='(-5e-3*mc_sig_vth-30e-3*mc_sig_vthp)*sw_stat_global*mc_skew'
.param pmos_3p3_sig_vth3='(-5e-3*mc_sig_vth-18e-3*mc_sig_vthp)*sw_stat_global*mc_skew'
.param pmos_3p3_tox='7.9e-009+(1.6e-10*mc_toxe+0.3e-10*mc_toxep)*sw_stat_global*mc_skew'
.param pmos_3p3_xl='(7e-9*mc_xl+4e-9*mc_xlp)*sw_stat_global*mc_skew'
.param pmos_3p3_xw='(7e-9*mc_xw+3e-9*mc_xwp)*sw_stat_global*mc_skew'
.param pmos_3p3_xj='1.0e-7+(0.3e-9*mc_xj+0.7e-9*mc_xjp)*sw_stat_global*mc_skew'
.param pmos_3p3_rdsw='466*(1+0.15*mc_rdswp*sw_stat_global*mc_skew)'
.param pmos_3p3_vth0_0='-0.7506174+pmos_3p3_sig_vth1'
.param pmos_3p3_vth0_1='-0.78216327+pmos_3p3_sig_vth1'
.param pmos_3p3_vth0_2='-0.76745877+pmos_3p3_sig_vth2'
.param pmos_3p3_vth0_3='-0.76841429+pmos_3p3_sig_vth2'
.param pmos_3p3_vth0_4='-0.7710094+pmos_3p3_sig_vth1'
.param pmos_3p3_vth0_5='-0.77464237+pmos_3p3_sig_vth2'
.param pmos_3p3_vth0_6='-0.77376777+pmos_3p3_sig_vth2'
.param pmos_3p3_vth0_7='-0.77390514+pmos_3p3_sig_vth3'
.param pmos_3p3_vth0_8='-0.76226585+pmos_3p3_sig_vth2'
.param pmos_3p3_vth0_9='-0.76552347+pmos_3p3_sig_vth2'
.param pmos_3p3_vth0_10='-0.7677531+pmos_3p3_sig_vth3'
.param pmos_3p3_vth0_11='-0.7682+pmos_3p3_sig_vth3'
.param pmos_3p3_vth0_12='-0.76184364+pmos_3p3_sig_vth2'
.param pmos_3p3_vth0_13='-0.76642857+pmos_3p3_sig_vth3'
.param pmos_3p3_vth0_14='-0.76779091+pmos_3p3_sig_vth3'
.param pmos_3p3_vth0_15='-0.7682+pmos_3p3_sig_vth3'
.param nmos_6p0_vsat='(1-0.063*mc_rdswn*sw_stat_global*mc_skew)'
.param nmos_6p0_vth0='(8e-3*mc_sig_vth+28e-3*mc_sig_vthn)*sw_stat_global*mc_skew'
.param nmos_6p0_xl='(2e-8*mc_xl+0*mc_xln)*sw_stat_global*mc_skew'
.param nmos_6p0_xw='(1.5e-8*mc_xw+9e-9*mc_xwn)*sw_stat_global*mc_skew'
.param nmos_6p0_tox='(4e-10*mc_toxe+1.3e-10*mc_toxen)*sw_stat_global*mc_skew'
.param nmos_6p0_cgso=1
.param nmos_6p0_cgdo=1
.param pmos_6p0_vth0='-0.8978+(8e-3*mc_sig_vth+30e-3*mc_sig_vthp)*sw_stat_global*mc_skew'
.param pmos_6p0_tox='156e-010+(4e-10*mc_toxe+1e-10*mc_toxep)*sw_stat_global*mc_skew'
.param pmos_6p0_xl='0+(2e-8*mc_xl+2e-9*mc_xlp)*sw_stat_global*mc_skew'
.param pmos_6p0_xw='0+(1.5e-8*mc_xw+9e-9*mc_xwp)*sw_stat_global*mc_skew'
.param pmos_6p0_xj='1.5e-7+(0.3e-9*mc_xj+1e-8*mc_xjp)*sw_stat_global*mc_skew'
.param pmos_6p0_rdsw='1426*(1+0.2*mc_rdswp*sw_stat_global*mc_skew)'
.param nmos_6p0_nat_vth0='-0.039+(8e-3*mc_sig_vth+60e-3*mc_sig_vthn)*sw_stat_global*mc_skew'
.param nmos_6p0_nat_tox='152e-010+(4e-10*mc_toxe+6e-10*mc_toxen)*sw_stat_global*mc_skew'
.param nmos_6p0_nat_xl='0+(2e-8*mc_xl+8e-8*mc_xln)*sw_stat_global*mc_skew'
.param nmos_6p0_nat_xw='0+(1.5e-8*mc_xw+8e-8*mc_xwn)*sw_stat_global*mc_skew'
.param nmos_6p0_nat_xj='1.5e-7+(0.3e-9*mc_xj+2e-8*mc_xjn)*sw_stat_global*mc_skew'
.param nmos_6p0_nat_rdsw='3480*(1+0.2*mc_rdswn*sw_stat_global*mc_skew)'
.param rsh_nplus2_u=60
.param rsh_pplus2_u=185
.param rsh_nplus_u_m='rsh_nplus2_u*(1+(mc_rsh_nplus_u/(rsh_nplus2_u))*res_mc_skew*sw_stat_global)'
.param rsh_pplus_u_m='rsh_pplus2_u*(1+(mc_rsh_pplus_u/(rsh_pplus2_u))*res_mc_skew*sw_stat_global)'
.lib 'sm141064.spice' fets_mm
.lib 'sm141064.spice' nmos_3p3_stat
.lib 'sm141064.spice' pmos_3p3_stat
.lib 'sm141064.spice' nmos_6p0_t
.lib 'sm141064.spice' pmos_6p0_stat
.lib 'sm141064.spice' nmos_6p0_nat_stat
.lib 'sm141064.spice' noise_corner
.endl statistical

.lib noise_corner
.param nmos_3p3_noia='(fnoicor==0)*3.2e+041+(fnoicor==1)*3.5e+042'
.param nmos_3p3_noib='(fnoicor==0)*1.2e+020+(fnoicor==1)*1.2e+020'
.param nmos_3p3_noic='(fnoicor==0)*6.0e+008+(fnoicor==1)*6.0e+008'
.param pmos_3p3_noia='(fnoicor==0)*3.2e+041+(fnoicor==1)*4.0e+042'
.param pmos_3p3_noib='(fnoicor==0)*1.8e+020+(fnoicor==1)*1.8e+020'
.param pmos_3p3_noic='(fnoicor==0)*3.0e+009+(fnoicor==1)*6.0e+009'
.param nmos_6p0_noia='(fnoicor==0)*1.998e+041+(fnoicor==1)*8e+041'
.param nmos_6p0_noib='(fnoicor==0)*1e+025+(fnoicor==1)*4e+025'
.param nmos_6p0_noic='(fnoicor==0)*5e+008+(fnoicor==1)*2e+009'
.param pmos_6p0_noia='(fnoicor==0)*6e+040+(fnoicor==1)*2e+043'
.param pmos_6p0_noib='(fnoicor==0)*1.5945e+025+(fnoicor==1)*1.5945e+025'
.param pmos_6p0_noic='(fnoicor==0)*1.0499e+009+(fnoicor==1)*1.0499e+009'
.param nmos_6p0_nat_noia='(fnoicor==0)*5.5e+040+(fnoicor==1)*1e+041'
.param nmos_6p0_nat_noib='(fnoicor==0)*2.5e+025+(fnoicor==1)*9.5e+025'
.param nmos_6p0_nat_noic='(fnoicor==0)*1e+007+(fnoicor==1)*2e+007'
.endl noise_corner

.lib nmos_3p3_t
.subckt nmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.007148
.param par_k=0.007008
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b nplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b nplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b nmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model nmos_3p3.0 nmos a0=0.11197377 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.32403844 alpha0=2.652013e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=19.905584 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0036363636 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95938091 k2=0.054714558 k3=0 k3b=0 keta=-0.14896036 kt1=-0.45934558 kt1l=0 kt2=-0.024730519 ku0=0 kvsat=0 kvth0=0 la0=-3.1454545e-009 lags=-1.5116364e-008 lalpha0=-3.0506364e-013 lbeta0=1.2863636e-007 ldelta=3.1818182e-009 level=54 lint=0 lk1=-9.9985454e-008 lk2=-4.1647636e-008 lketa=3.8830182e-008 lkt1=4.2126364e-008 lkt2=1.2545455e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-4.729e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.6525455e-009 lua=7.0220545e-016 lub1=2.8745455e-025 lub=-7.9058636e-025 luc1=-3.8181818e-018 luc=-6.1360545e-017 lute=9.0909091e-008 lvoff=3.9354545e-009 lvsat=-0.0027272727 lvth0=-3.8715455e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.7450182e-015 pags=-1.2213818e-014 palpha0=-1.3658182e-020 paramchk=1 pbeta0=8.7272727e-016 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.3741 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=5.388e-015 pketa=-2.4261818e-015 pkt1=-8.6530909e-015 pkt2=-2.9672727e-016 ppclm=8.5658182e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-6.5127273e-016 pua=-1.4149745e-022 pub1=-5.7490909e-032 pub=9.2644364e-032 puc1=1.8327273e-024 puc=5.4467782e-024 pute=-4.3636364e-014 pvag=0 pvoff=-1.4858182e-015 pvsat=1.3090909e-009 pvth0=4.3636364e-016 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.023671338 ua1=1.675e-009 ua=-1.1554452e-009 ub1=-4.1945234e-018 ub=3.3771156e-018 uc1=-4.2363636e-011 uc=2.2660166e-010 ute=-1.5675325 vbm=-3 version=4.5 vfbcv=-1 voff=-0.1262652 voffcv=0.005 voffl=0 vsat=92454.546 vth0=0.70837662 w0=5e-007 wa0=-6.2322078e-009 wags=4.7930493e-008 walpha0=4.8779221e-014 wbeta0=1.3848312e-007 wint=1e-008 wk2=-1.9242857e-008 wketa=8.1643636e-009 wkt1=3.2086753e-008 wkt2=1.0597403e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.1028364e-008 wr=1 wtvoff=0 wu0=4.6066597e-009 wua=2.7073777e-016 wub1=3.3492467e-025 wub=-4.093733e-025 wuc1=-6.5454545e-018 wuc=-3.2577351e-017 wute=1.0441558e-007 wvoff=5.3064935e-009 wvsat=-0.00021818182 wvth0=-1.430587e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.1 nmos a0=1.0861147 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.47870122 alpha0=6.5720816e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=22.625306 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0014285714 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.74639857 k2=0.0237458 k3=0 k3b=0 keta=-0.028417143 kt1=-0.33916633 kt1l=0 kt2=-0.020311225 ku0=0 kvsat=0 kvth0=0 la0=-4.9021592e-007 lags=-9.2447755e-008 lalpha0=-2.265098e-012 lbeta0=-1.2312245e-006 ldelta=4.2857143e-009 level=54 lint=0 lk1=6.5057143e-009 lk2=-2.6163257e-008 lketa=-2.1441429e-008 lkt1=-1.7963265e-008 lkt2=-9.5510204e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=9.8313061e-008 lpdiblc2=9.06e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.6503673e-009 lua=7.7258204e-016 lub1=-4.0760816e-025 lub=-6.4387347e-025 luc1=5.1428571e-018 luc=9.6333061e-018 lvoff=-2.8273469e-009 lvsat=0.0017142857 lvth0=-2.3433061e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.4627526e-014 pags=-9.9007347e-015 palpha0=1.8396735e-020 paramchk=1 pbeta0=2.4538775e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.082893878 pdiblc1=0.39 pdiblc2=0.001359 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=-2.7269486e-015 pketa=5.3691429e-015 pkt1=8.6223674e-015 pkt2=2.5273469e-016 ppclm=-2.8711837e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.2234122e-015 pua=-2.976098e-023 pub1=8.1521633e-032 pub=-9.8501878e-032 puc1=-2.4685714e-024 puc=-1.1961815e-023 pvag=0 pvoff=3.2032653e-016 pvsat=2.0571429e-009 pvth0=-5.642449e-016 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.029675694 ua1=1.675e-009 ua=-1.2961984e-009 ub1=-2.804398e-018 ub=3.0836898e-018 uc1=-6.0285714e-011 uc=8.4613959e-011 ute=-1.3857143 vbm=-3 version=4.5 vfbcv=-1 voff=-0.11273959 voffcv=0.005 voffl=0 vsat=83571.429 vth0=0.67781184 w0=5e-007 wa0=-5.1997224e-008 wags=4.3304327e-008 walpha0=-1.5330612e-014 wbeta0=-3.5054694e-007 wint=1e-008 wk2=-3.01296e-009 wketa=-7.4262857e-009 wkt1=-2.4641633e-009 wkt2=-3.9183673e-011 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=4.3902367e-008 wr=1 wtvoff=0 wu0=8.572898e-010 wua=4.7264816e-017 wub1=5.6899592e-026 wub=-2.7080816e-026 wuc1=2.0571429e-018 wuc=2.2398367e-018 wute=1.7142857e-008 wvoff=1.6942041e-009 wvsat=-0.0017142857 wvth0=-1.2304653e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.2 nmos a0=1.224418 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.25784649 alpha0=7.5243347e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.210162 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027272727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79593364 k2=0.0056393844 k3=0 k3b=0 keta=-0.019651071 kt1=-0.32898149 kt1l=0 kt2=-0.021107143 ku0=0 kvsat=0 kvth0=0 la0=-6.5617987e-007 lags=1.7257792e-007 lalpha0=-8.4670617e-011 lbeta0=-3.133052e-006 ldelta=2.7272727e-009 level=54 lint=0 lk1=-5.2936364e-008 lk2=-4.4355584e-009 lketa=-3.1960714e-008 lkt1=-3.0185065e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=-2.9236364e-008 lpdiblc2=1.7686364e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.6755195e-009 lua=1.9570909e-016 lub1=-7.5296104e-025 lub=-2.347987e-025 luc=-6.9921429e-018 lvoff=1.3461039e-008 lvth0=-3.224026e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-4.2919481e-014 pags=4.5191688e-014 palpha0=-9.043013e-018 paramchk=1 pbeta0=-3.1184416e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.18918506 pdiblc1=0.39 pdiblc2=0.00064013636 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=2.6091117e-015 pketa=-2.7504935e-015 pkt1=1.4488831e-014 ppclm=4.7225454e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.447013e-015 pua=1.9701818e-023 pub1=1.231013e-031 pub=-1.1174026e-031 puc=1.4030649e-024 pvag=0 pvoff=-1.4493507e-016 pvth0=-3.6888312e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032447266 ua1=1.675e-009 ua=-8.1547091e-010 ub1=-2.5166039e-018 ub=2.7427942e-018 uc1=-5.6e-011 uc=9.84685e-011 ute=-1.3857143 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12631325 voffcv=0.005 voffl=0 vsat=85000 vth0=0.66097097 w0=5e-007 wa0=4.291948e-009 wags=-2.606026e-009 walpha0=7.5358442e-012 wbeta0=1.1381299e-007 wint=1e-008 wk2=-7.4596769e-009 wketa=-6.5992208e-010 wkt1=-7.3528831e-009 wkt2=1.7142857e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.1551688e-009 wr=1 wtvoff=0 wu0=6.7095584e-010 wua=6.0458182e-018 wub1=2.224987e-026 wub=-1.6048831e-026 wuc=-8.8975636e-018 wute=1.7142857e-008 wvoff=2.0819221e-009 wvth0=-9.7008312e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.3 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.27510429 alpha0=6.6776286e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.896857 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=0.0051958286 k3=0 k3b=0 keta=-0.022847143 kt1=-0.332 kt1l=0 kt2=-0.021107143 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.18626143 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032279714 ua1=1.675e-009 ua=-7.959e-010 ub1=-2.5919e-018 ub=2.7193143e-018 uc1=-5.6e-011 uc=9.7769286e-011 ute=-1.3857143 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12496714 voffcv=0.005 voffl=0 vsat=85000 vth0=0.66064857 w0=5e-007 wags=1.9131429e-009 walpha0=6.6315429e-012 wbeta0=8.2628571e-008 wint=1e-008 wk2=-7.1987657e-009 wketa=-9.3497143e-010 wkt1=-5.904e-009 wkt2=1.7142857e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=6.8777143e-009 wr=1 wtvoff=0 wu0=8.1565714e-010 wua=8.016e-018 wub1=3.456e-026 wub=-2.7222857e-026 wuc=-8.7572571e-018 wute=1.7142857e-008 wvoff=2.0674286e-009 wvth0=-1.0069714e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.4 nmos a0=0.10680558 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.35500309 alpha0=2.6500109e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=20.982852 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0036363636 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95938091 k2=0.041255727 k3=0 k3b=0 keta=-0.12490989 kt1=-0.37773746 kt1l=0 kt2=-0.014603854 ku0=0 kvsat=0 kvth0=0 la0=-1.6983636e-009 lags=-1.1780546e-008 lalpha0=-2.8170545e-013 lbeta0=-8.9454546e-008 ldelta=3.1818182e-009 level=54 lint=0 lk1=-9.9985454e-008 lk2=-3.7879164e-008 lketa=3.0254945e-008 lkt1=1.6718727e-008 lkt2=-3.3230727e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-8.0088e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.0251818e-009 lua=3.9938436e-016 lub1=2.4878e-025 lub=-9.0230909e-026 luc=-3.4349127e-017 lvoff=-9.2114546e-009 lvsat=0.0042909091 lvth0=-4.1979273e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.0504145e-015 pags=-1.3815011e-014 palpha0=-2.4870109e-020 paramchk=1 pbeta0=1.0555636e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.45921829 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=3.5791331e-015 pketa=1.6899316e-015 pkt1=3.5425745e-015 pkt2=1.9005294e-015 ppclm=2.4308858e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.5013818e-016 pua=3.8566691e-024 pub1=-3.8927127e-032 pub=-2.4352626e-031 puc=-7.5187026e-024 pvag=0 pvoff=4.8246982e-015 pvsat=-2.0596364e-009 pvth0=2.0029964e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.033011551 ua1=1.675e-009 ua=-6.3005701e-010 ub1=-3.65896e-018 ub=2.2836418e-018 uc1=-5.6e-011 uc=1.5877203e-010 ute=-1.4342857 vbm=-3 version=4.5 vfbcv=-1 voff=-0.079311948 voffcv=0.005 voffl=0 vsat=71618.182 vth0=0.72356597 w0=5e-007 wa0=-3.7514805e-009 wags=3.3067462e-008 walpha0=4.9740218e-014 wbeta0=-3.786053e-007 wint=1e-008 wk2=-1.2782618e-008 wketa=-3.3798633e-009 wkt1=-7.0851491e-009 wkt2=-3.8010589e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.9828414e-008 wr=1 wtvoff=0 wu0=1.2335751e-010 wua=1.8551439e-017 wub1=7.7854254e-026 wub=1.1549411e-025 wuc=-1.9125195e-020 wute=4.0457143e-008 wvoff=-1.7231065e-008 wvsat=0.0097832727 wvth0=-2.1596758e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.5 nmos a0=0.97533082 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.441074 alpha0=6.8164074e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.036008 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0014285714 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.76833212 k2=0.0082103273 k3=0 k3b=0 keta=-0.043888571 kt1=-0.4079911 kt1l=0 kt2=-0.031229592 ku0=0 kvsat=0 kvth0=0 la0=-4.3596098e-007 lags=-5.4816e-008 lalpha0=-2.3649037e-012 lbeta0=-1.1603265e-007 ldelta=4.2857143e-009 level=54 lint=0 lk1=-4.4610612e-009 lk2=-2.1356464e-008 lketa=-1.0255714e-008 lkt1=3.1845551e-008 lkt2=4.9897959e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=4.0921959e-008 lpdiblc2=9.06e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.9403755e-009 lua=6.6367861e-016 lub1=-1.7578531e-025 lub=-3.6042122e-025 luc1=3.1443869e-017 luc=4.0383673e-018 lvoff=1.1378694e-008 lvsat=-0.0041142857 lvth0=-1.7716408e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.4148441e-015 pags=-2.7963977e-014 palpha0=6.6303478e-020 paramchk=1 pbeta0=-2.8990433e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21719837 pdiblc1=0.39 pdiblc2=0.001359 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=5.2640522e-015 pk2=-5.0342094e-015 pkt1=-1.5285865e-014 pkt2=-2.6008163e-015 ppclm=2.4676545e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.5579167e-016 pua=2.2512666e-023 pub1=-2.9753339e-032 pub=-2.3455895e-031 puc1=-1.5093057e-023 puc=-9.2762449e-024 pvag=0 pvoff=-6.4985731e-015 pvsat=4.8548571e-009 pvth0=-3.3082384e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.031181163 ua1=1.675e-009 ua=-1.1586455e-009 ub1=-2.8098294e-018 ub=2.8240225e-018 uc1=-1.1888774e-010 uc=8.1997037e-011 ute=-1.4342857 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12049225 voffcv=0.005 voffl=0 vsat=88428.571 vth0=0.67504024 w0=5e-007 wa0=1.1790367e-009 wags=6.1365394e-008 walpha0=-1.3260696e-013 wbeta0=4.1231608e-007 wint=1e-008 wk1=-1.0528104e-008 wk2=4.4440669e-009 wkt1=3.0571729e-008 wkt2=5.2016327e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-2.0563788e-008 wr=1 wtvoff=0 wu0=1.3466449e-010 wua=-1.8760555e-017 wub1=5.9506678e-026 wub=9.755951e-026 wuc1=3.0186115e-017 wuc=3.4959595e-018 wute=4.0457143e-008 wvoff=5.4154776e-009 wvsat=-0.0040457143 wvth0=-1.0974289e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.6 nmos a0=1.2333595 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.28370796 alpha0=9.0921047e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.039866 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027272727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79418892 k2=-0.0057236965 k3=0 k3b=0 keta=-0.021025909 kt1=-0.33923366 kt1l=0 kt2=-0.021803571 ku0=0 kvsat=0 kvth0=0 la0=-7.4559545e-007 lags=1.3402325e-007 lalpha0=-1.0329047e-010 lbeta0=-3.7206623e-006 ldelta=2.7272727e-009 level=54 lint=0 lk1=-3.5489221e-008 lk2=-4.6356351e-009 lketa=-3.7690909e-008 lkt1=-5.0663377e-008 lkt2=-6.3214286e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=2.9060649e-008 lpdiblc2=1.7686364e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.4308442e-009 lua=2.1903156e-016 lub1=7.0824935e-025 lub=-6.4298182e-025 luc1=-5.0024338e-017 luc=-1.4633922e-017 lute=3.448052e-007 lvoff=1.3159091e-008 lvth0=1.325026e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=6.3697932e-014 palpha0=-1.0548281e-019 paramchk=1 pbeta0=-2.9791169e-014 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.22708279 pdiblc1=0.39 pdiblc2=0.00064013636 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-8.3746286e-015 pk2=2.7051485e-015 pkt1=2.4318421e-014 pkt2=3.0342857e-015 ppclm=1.9242888e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.3295688e-015 pua=8.5070338e-024 pub1=-5.7827969e-031 pub=8.4187636e-032 puc1=2.4011682e-023 puc=5.071119e-024 pute=-1.6550649e-013 pvag=0 pvth0=-1.1596488e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.036490513 ua1=1.675e-009 ua=-7.881063e-010 ub1=-3.5465249e-018 ub=3.0594896e-018 uc1=-5.0997566e-011 uc=9.7557278e-011 ute=-1.7216234 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12197591 voffcv=0.005 voffl=0 vsat=85000 vth0=0.64923469 w0=5e-007 wags=-1.501953e-008 walpha0=1.0548281e-014 wbeta0=1.9555512e-007 wint=1e-008 wk1=8.3746286e-010 wk2=-2.005398e-009 wkt1=-2.4318421e-009 wkt2=5.0571429e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.603574e-008 wr=1 wtvoff=0 wu0=-1.2698026e-009 wua=-7.0891948e-018 wub1=5.1661197e-025 wub=-1.6806265e-025 wuc1=-2.4011682e-018 wuc=-8.460177e-018 wute=1.7837922e-007 wvth0=-4.067414e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.7 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29711029 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.6678 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=-0.00618726 k3=0 k3b=0 keta=-0.024795 kt1=-0.3443 kt1l=0 kt2=-0.022435714 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.22998886 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.036347429 ua1=1.675e-009 ua=-7.6620314e-010 ub1=-3.4757e-018 ub=2.9951914e-018 uc1=-5.6e-011 uc=9.6093886e-011 ute=-1.6871429 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.005 voffl=0 vsat=85000 vth0=0.65055971 w0=5e-007 wags=-8.6497371e-009 wbeta0=1.92576e-007 wint=1e-008 wk2=-1.7348832e-009 wkt2=8.0914286e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.4111451e-008 wr=1 wtvoff=0 wu0=-1.1368457e-009 wua=-6.2384914e-018 wub1=4.58784e-025 wub=-1.5964389e-025 wuc=-7.9530651e-018 wute=1.6182857e-007 wvth0=-5.2270629e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.8 nmos a0=0.10362636 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.2705431 alpha0=2.5953123e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.140586 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0036363636 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95060511 k2=0.013945175 k3=0 k3b=0 keta=-0.12424077 kt1=-0.28115299 kt1l=0 kt2=-0.025449687 ku0=0 kvsat=0 kvth0=0 la0=-8.0818182e-010 lags=3.2753448e-008 lalpha0=-2.5435614e-013 ldelta=3.1818182e-009 level=54 lint=0 lk1=-9.5597554e-008 lk2=-3.0232209e-008 lketa=2.9920384e-008 lkt1=-1.0099496e-008 lkt2=9.6575269e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.2990496e-006 lpclm=-9.798626e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.7050207e-010 lua=2.5458994e-016 lub1=4.827456e-025 lub=-3.3240512e-025 luc1=4.973267e-017 luc=-6.8059408e-017 lvoff=6.8691116e-010 lvoffcv=-1.118626e-007 lvsat=-0.00034132231 lvth0=-5.5747725e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.59809917 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=-6.6365124e-014 palpha0=-5.7142305e-020 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.20476889 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-5.177723e-015 pk2=-5.4442735e-015 pketa=2.0847148e-015 pkt1=3.5188078e-014 pkt2=-3.1602845e-015 pnoff=-1.5328785e-012 ppclm=-5.8632603e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=4.1983839e-015 pua=1.7471409e-022 pub1=-3.1500653e-031 pub=4.2239319e-032 puc1=-5.8684551e-023 puc=3.2259428e-023 pvag=0 pvoff=-6.8553733e-015 pvoffcv=1.3199787e-013 pvsat=3.4063967e-009 pvth0=1.824977e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.046898182 ua1=1.675e-009 ua=-6.6207759e-010 ub1=-5.3788142e-018 ub=3.7962141e-018 uc1=-2.2938539e-010 uc=2.9436835e-010 ute=-1.5701136 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12424632 voffcv=0.22872521 voffl=0 vsat=85682.645 vth0=0.75419347 w0=5e-007 wags=1.3273025e-007 walpha0=1.1428461e-013 wbeta0=-5.6473191e-007 wint=1e-008 wk1=1.0355446e-008 wk2=1.9443834e-008 wketa=-4.1694295e-009 wkt1=-1.2105482e-007 wkt2=8.9970236e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=3.065757e-006 wpclm=2.8042187e-007 wr=1 wtvoff=0 wu0=-1.6262868e-008 wua=5.6335718e-017 wub1=2.1072821e-024 wub=-1.6693412e-024 wuc1=2.0459475e-016 wuc=-1.6002278e-016 wute=2.0073409e-007 wvoff=3.5791497e-008 wvoffcv=-2.6399574e-007 wvsat=-0.0068127934 wvth0=-5.7737207e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.9 nmos a0=0.57970277 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.63340774 alpha0=6.7040286e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.043581 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0014285714 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.017155231 k3=0 k3b=0 keta=-0.043888571 kt1=-0.30297354 kt1l=0 kt2=-0.021799026 ku0=0 kvsat=0 kvth0=0 la0=-2.3884638e-007 lags=-1.4867887e-007 lalpha0=-2.3087143e-012 lbeta0=4.8502597e-008 ldelta=4.2857143e-009 level=54 lint=0 lk2=-3.1837237e-008 lketa=-1.0255714e-008 lkt1=8.1077922e-010 lkt2=-8.5957792e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=6.8726318e-008 lpdiblc2=9.06e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.387089e-009 lua=3.880134e-016 lub1=-6.899552e-025 lub=-1.7056325e-025 luc1=7.5986727e-018 luc=5.1261039e-019 lvoff=-1.0167857e-008 lvth0=-9.953513e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.3401007e-013 pags=8.279421e-014 paramchk=1 pbeta0=-4.8405592e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.047719 pdiblc1=0.39 pdiblc2=0.001359 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=7.3331031e-015 pkt1=2.1335166e-014 pkt2=4.3014448e-015 ppclm=-8.1325983e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=2.9708645e-016 pua=3.4779762e-022 pub1=5.7696713e-031 pub=-4.5859137e-031 puc1=1.3044275e-023 puc=-5.1158517e-024 pvag=0 pvoff=1.8926357e-014 pvth0=-1.2468455e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.038465008 ua1=1.675e-009 ua=-9.289245e-010 ub1=-3.0334126e-018 ub=3.4725304e-018 uc1=-1.4511739e-010 uc=1.5722431e-010 ute=-1.5701136 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10253679 voffcv=0.005 voffl=0 vsat=85000 vth0=0.66260505 w0=5e-007 wa0=4.6802014e-007 wags=-1.6558842e-007 wbeta0=4.0337993e-007 wint=1e-008 wk2=-6.1109193e-009 wkt1=-9.3348999e-008 wkt2=-5.9264351e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.7942187e-007 wr=1 wtvoff=0 wu0=-8.4602728e-009 wua=-2.8983135e-016 wub1=3.2333483e-025 wub=-6.6767982e-025 wuc1=6.1137104e-017 wuc=-8.5272224e-017 wute=2.0073409e-007 wvoff=-1.5771964e-008 wvth0=3.6992425e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.10 nmos a0=1.175342 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26729169 alpha0=9.0929986e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.512311 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027272727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79747612 k2=-0.0074231864 k3=0 k3b=0 keta=-0.021025909 kt1=-0.31506405 kt1l=0 kt2=-0.016812862 ku0=0 kvsat=0 kvth0=0 la0=-9.536135e-007 lags=2.9066039e-007 lalpha0=-1.0337986e-010 lbeta0=-4.1139731e-006 ldelta=2.7272727e-009 level=54 lint=0 lk1=-4.5679339e-008 lk2=-2.3431364e-009 lketa=-3.7690909e-008 lkt1=1.5319401e-008 lkt2=-6.8429752e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.5464876e-007 lpclm=-1.5414418e-007 lpdiblc2=1.7686364e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.9522345e-009 lua1=2.5980992e-017 lua=2.4617513e-016 lub1=-1.7520434e-024 lub=1.6897655e-025 luc1=-1.1288886e-016 luc=6.3987831e-017 lute=-2.7427686e-008 lvoff=1.3159091e-008 lvoffcv=8.5056818e-008 lvth0=7.3817355e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.128874 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.454613e-013 pags=-1.211339e-013 paramchk=1 pbeta0=4.3431558e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23344442 pdiblc1=0.39 pdiblc2=0.00064013636 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=3.6497107e-015 pkt1=-5.3541257e-014 pkt2=3.6497107e-015 pnoff=1.8248554e-013 ppclm=2.3542459e-013 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-2.662464e-015 pua1=-3.065757e-023 pua=-2.3522386e-023 pub1=2.3248657e-030 pub=-8.7392324e-031 puc1=9.8191818e-023 puc=-8.7702549e-023 pute=2.7372831e-013 pvag=0 pvoffcv=-1.0036705e-013 pvth0=-4.6716298e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040494054 ua1=1.6533492e-009 ua=-8.1072595e-010 ub1=-2.1483391e-018 ub=3.1895805e-018 uc1=-4.4711114e-011 uc=1.0432829e-010 ute=-1.5472572 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12197591 voffcv=-0.065880682 voffl=0 vsat=85000 vth0=0.64815901 w0=5e-007 wa0=6.8460666e-008 wags=4.3516718e-009 wbeta0=-3.6192965e-007 wint=1e-008 wk1=-3.0414256e-009 wkt1=-3.095198e-008 wkt2=-5.3833233e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.5207128e-007 wpclm=-2.3542459e-008 wr=1 wtvoff=0 wu0=-5.9939808e-009 wua1=2.5547975e-017 wua=1.9601988e-017 wub1=-1.1332474e-024 wub=-3.2156993e-025 wuc1=-9.8191818e-018 wuc=-1.6449976e-017 wute=-2.7372831e-008 wvoffcv=8.3639205e-008 wvth0=-2.7981116e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.11 nmos a0=1.0799807 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29635773 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.100914 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79290818 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31353211 kt1l=0 kt2=-0.017497159 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1134091 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040689277 ua1=1.6559473e-009 ua=-7.8610843e-010 ub1=-2.3235434e-018 ub=3.2064782e-018 uc1=-5.6e-011 uc=1.1072708e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.057375 voffl=0 vsat=85000 vth0=0.64889718 w0=5e-007 wa0=9.3006796e-008 wags=-7.7617182e-009 wbeta0=-3.1849809e-007 wint=1e-008 wk1=-2.6764545e-009 wkt1=-3.6306106e-008 wkt2=-5.0183523e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.3382273e-007 wr=1 wtvoff=0 wu0=-6.2602272e-009 wua1=2.2482218e-017 wua=1.7249749e-017 wub1=-9.0076078e-025 wub=-4.0896225e-025 wuc=-2.5220231e-017 wvoffcv=7.36025e-008 wvth0=-3.2652745e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.12 nmos a0=0.13211844 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.46155061 alpha0=2.6067636e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=2.3e-010 cgidl=0.5 cgsl=1e-010 cgso=2.3e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0036363636 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95164273 k2=0.015893454 k3=0 k3b=0 keta=-0.12105603 kt1=-0.29328273 kt1l=0 kt2=-0.024548182 ku0=0 kvsat=0 kvth0=0 la0=-1.5054221e-008 lags=-6.2750307e-008 lalpha0=-2.6008182e-013 ldelta=3.1818182e-009 level=54 lint=0 lk1=-9.6116364e-008 lk2=-3.0777727e-008 lketa=2.8328017e-008 lkt1=-6.5736364e-009 lkt2=6.4909091e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.1454545e-006 lpclm=-1.5673636e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=5.9118182e-010 lua=2.7209636e-016 lub1=4.5118182e-025 lub=-3.2817273e-025 luc1=4.3852454e-017 luc=-6.4827e-017 lvoffcv=-9.8636364e-008 lvth0=-5.3919091e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.29090909 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.4217547e-013 pags=8.8676235e-013 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23286727 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pketa=1.7976533e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.045268636 ua1=1.675e-009 ua=-6.5643273e-010 ub1=-5.1676636e-018 ub=3.6289455e-018 uc1=-2.0888491e-010 uc=2.78334e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.20227273 voffl=0 vsat=85000 vth0=0.74840818 w0=5e-007 wa0=-2.8435094e-007 wags=-1.7735247e-006 wint=1e-008 wketa=-3.5953066e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.13 nmos a0=0.62659857 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.61681571 alpha0=6.7040286e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0014285714 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.016542914 k3=0 k3b=0 keta=-0.043888571 kt1=-0.31232714 kt1l=0 kt2=-0.022392857 ku0=0 kvsat=0 kvth0=0 la0=-2.6229429e-007 lags=-1.4038286e-007 lalpha0=-2.3087143e-012 ldelta=4.2857143e-009 level=54 lint=0 lk2=-3.1102457e-008 lketa=-1.0255714e-008 lkt1=2.9485714e-009 lkt2=-4.2857143e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=6.7911429e-008 lpdiblc2=9.06e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.4168571e-009 lua=4.2286286e-016 lub1=-6.3214286e-025 lub=-2.1651429e-025 luc1=8.9057143e-018 lvoff=-8.2714286e-009 lvth0=-1.1202857e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.065697143 pdiblc1=0.39 pdiblc2=0.001359 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.037617286 ua1=1.675e-009 ua=-9.5796571e-010 ub1=-3.0010143e-018 ub=3.4056286e-018 uc1=-1.3899143e-010 uc=1.4868e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10411714 voffcv=0.005 voffl=0 vsat=85000 vth0=0.66297571 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.14 nmos a0=1.1822018 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26772773 alpha0=9.0929986e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.476046 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027272727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79717136 k2=-0.0074231864 k3=0 k3b=0 keta=-0.021025909 kt1=-0.31816545 kt1l=0 kt2=-0.017352273 ku0=0 kvsat=0 kvth0=0 la0=-9.2901818e-007 lags=2.7852273e-007 lalpha0=-1.0337986e-010 lbeta0=-4.0704545e-006 ldelta=2.7272727e-009 level=54 lint=0 lk1=-4.5313636e-008 lk2=-2.3431364e-009 lketa=-3.7690909e-008 lkt1=9.9545454e-009 lkt2=-6.4772727e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.3636364e-007 lpclm=-1.3055455e-007 lpdiblc2=1.7686364e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.6854546e-009 lua1=2.2909091e-017 lua=2.4381818e-016 lub1=-1.5190909e-024 lub=8.1409091e-026 luc1=-1.0305e-016 luc=5.52e-017 lvoff=1.3159091e-008 lvoffcv=7.5e-008 lvth0=6.9136364e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1136364 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23108545 pdiblc1=0.39 pdiblc2=0.00064013636 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.039893455 ua1=1.6559091e-009 ua=-8.0876182e-010 ub1=-2.2618909e-018 ub=3.1573591e-018 uc1=-4.5695e-011 uc=1.0268e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12197591 voffcv=-0.0575 voffl=0 vsat=85000 vth0=0.64787864 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model nmos_3p3.15 nmos a0=1.0893 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29558 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.069 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=2.3e-010 cgidl=0.5 cgsl=1e-010 cgso=2.3e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79264 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31717 kt1l=0 kt2=-0.018 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8e-009 toxm=8e-009 toxp=8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040062 ua1=1.6582e-009 ua=-7.8438e-010 ub1=-2.4138e-018 ub=3.1655e-018 uc1=-5.6e-011 uc=1.082e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.05 voffl=0 vsat=85000 vth0=0.64857 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.subckt nplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 r_rsh0='rsh_nplus_u_m' r_dw=-5e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.36e-3 r_tc2=6.5e-7 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model np_junction d cj=0.00096797 level=2
d1 3 1 np_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends nplus_u_m1
.endl nmos_3p3_t

.lib nmos_3p3_f
.subckt nmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.007148
.param par_k=0.007008
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b nplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b nplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b nmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model nmos_3p3.0 nmos a0=0.11226647 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.31756239 alpha0=2.6143989e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=19.904932 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0039772727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.94866818 k2=0.052196642 k3=0 k3b=0 keta=-0.14562336 kt1=-0.45807784 kt1l=0 kt2=-0.024703182 ku0=0 kvsat=0 kvth0=0 la0=-3.0545135e-009 lags=-1.270937e-008 lalpha0=-2.787532e-013 lbeta0=1.1800932e-007 ldelta=2.9210227e-009 level=54 lint=0 lk1=-9.1790218e-008 lk2=-3.8749265e-008 lketa=3.5879506e-008 lkt1=3.950099e-008 lkt2=1.1800932e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-4.4233047e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.3334833e-009 lua=6.5818091e-016 lub1=2.6939132e-025 lub=-7.3464598e-025 luc1=-3.6804886e-018 luc=-5.6852041e-017 lute=8.7630682e-008 lvoff=3.7549747e-009 lvsat=-0.0026289205 lvth0=-3.5583899e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.717132e-015 pags=-1.2018636e-014 palpha0=-1.3439918e-020 paramchk=1 pbeta0=8.5878068e-016 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.36674716 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=5.3018972e-015 pketa=-2.3874103e-015 pkt1=-8.5148105e-015 pkt2=-2.9198543e-016 ppclm=8.4289324e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-6.4086508e-016 pua=-1.3923626e-022 pub1=-5.6572177e-032 pub=9.1163863e-032 puc1=1.8034394e-024 puc=5.3597361e-024 pute=-4.2939034e-014 pvag=0 pvoff=-1.4620741e-015 pvsat=1.288171e-009 pvth0=4.2939034e-016 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.023697233 ua1=1.675e-009 ua=-1.1068315e-009 ub1=-4.197971e-018 ub=3.334019e-018 uc1=-4.2111364e-011 uc=2.2336e-010 ute=-1.5681818 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12637972 voffcv=0.005 voffl=0 vsat=99670.454 vth0=0.63571386 w0=5e-007 wa0=-6.4797433e-009 wags=4.9972817e-008 walpha0=5.071667e-014 wbeta0=1.4853682e-007 wint=1e-008 wk2=-2.0007159e-008 wketa=8.4725454e-009 wkt1=3.3399235e-008 wkt2=1.1018318e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.3523508e-008 wr=1 wtvoff=0 wu0=4.8629688e-009 wua=2.7394695e-016 wub1=3.5239491e-025 wub=-4.2815738e-025 wuc1=-6.8054318e-018 wuc=-3.4293319e-017 wute=1.0690909e-007 wvoff=5.5172608e-009 wvsat=-8.3522727e-005 wvth0=-1.5283991e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.1 nmos a0=1.0792115 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.47190495 alpha0=6.5170032e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=22.630402 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0015357143 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.74656121 k2=0.02341267 k3=0 k3b=0 keta=-0.028193589 kt1=-0.33938118 kt1l=0 kt2=-0.020331679 ku0=0 kvsat=0 kvth0=0 la0=-4.7202287e-007 lags=-8.7565511e-008 lalpha0=-2.1715163e-012 lbeta0=-1.2038436e-006 ldelta=4.1051786e-009 level=54 lint=0 lk1=6.2316611e-009 lk2=-2.4789039e-008 lketa=-2.1073934e-008 lkt1=-1.8066891e-008 lkt2=-9.4008589e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=9.4458106e-008 lpdiblc2=8.6783475e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.4587752e-009 lua=7.4300653e-016 lub1=-3.9857179e-025 lub=-6.0692192e-025 luc1=5.172525e-018 luc=1.0421037e-017 lvoff=-2.7402067e-009 lvsat=0.0014368125 lvth0=-2.2389644e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.528563e-014 pags=-1.0165305e-014 palpha0=1.8888337e-020 paramchk=1 pbeta0=2.5194507e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.080786018 pdiblc1=0.39 pdiblc2=0.00138165 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=-2.7998188e-015 pketa=5.5126185e-015 pkt1=8.8527765e-015 pkt2=2.5948834e-016 ppclm=-2.9479082e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.2561046e-015 pua=-3.055626e-023 pub1=8.3700075e-032 pub=-1.0113407e-031 puc1=-2.5345373e-024 puc=-1.2281462e-023 pvag=0 pvoff=3.2888638e-016 pvsat=2.1121144e-009 pvth0=-5.793228e-016 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.029624466 ua1=1.675e-009 ua=-1.2817297e-009 ub1=-2.8207275e-018 ub=3.0706704e-018 uc1=-6.0365e-011 uc=8.4652626e-011 ute=-1.3875 vbm=-3 version=4.5 vfbcv=-1 voff=-0.11298759 voffcv=0.005 voffl=0 vsat=91287.5 vth0=0.60850921 w0=5e-007 wa0=-5.5074584e-008 wags=4.6151516e-008 walpha0=-1.5939525e-014 wbeta0=-3.6916688e-007 wint=1e-008 wk2=-3.3025902e-009 wketa=-7.8161737e-009 wkt1=-2.4102225e-009 wkt2=-3.52275e-011 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=4.6980911e-008 wr=1 wtvoff=0 wu0=9.5169113e-010 wua=4.9864474e-017 wub1=6.3173775e-026 wub=-3.1666793e-026 wuc1=2.13885e-018 wuc=2.0802857e-018 wute=1.8375e-008 wvoff=1.8245588e-009 wvsat=-0.001782375 wvth0=-1.320417e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.2 nmos a0=1.2231563 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.25832779 alpha0=7.4353703e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.194431 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027306818 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79586747 k2=0.0064105499 k3=0 k3b=0 keta=-0.019621922 kt1=-0.32825519 kt1l=0 kt2=-0.021125 ku0=0 kvsat=0 kvth0=0 la0=-6.4259738e-007 lags=1.6552342e-007 lalpha0=-8.2558005e-011 lbeta0=-3.0572184e-006 ldelta=2.689142e-009 level=54 lint=0 lk1=-5.2196247e-008 lk2=-4.6415264e-009 lketa=-3.123136e-008 lkt1=-3.1251192e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=-3.3678143e-008 lpdiblc2=1.7439086e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.8007167e-009 lua=1.9094925e-016 lub1=-7.5507747e-025 lub=-2.2003905e-025 luc=-7.0384932e-018 lvoff=1.3287723e-008 lvth0=-2.8000692e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-4.536112e-014 pags=4.7762591e-014 palpha0=-9.5574596e-018 paramchk=1 pbeta0=-3.2958461e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.18891787 pdiblc1=0.39 pdiblc2=0.00064234716 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=2.757541e-015 pketa=-2.9069659e-015 pkt1=1.5313084e-014 ppclm=4.9912056e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.5293319e-015 pua=2.0822632e-023 pub1=1.3010439e-031 pub=-1.1809703e-031 puc=1.4828837e-024 pvag=0 pvoff=-1.5318025e-016 pvth0=-3.8986845e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032375092 ua1=1.675e-009 ua=-8.1585861e-010 ub1=-2.5198788e-018 ub=2.744187e-018 uc1=-5.6e-011 uc=9.9386407e-011 ute=-1.3875 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12651327 voffcv=0.005 voffl=0 vsat=92500 vth0=0.59197793 w0=5e-007 wa0=4.5429264e-009 wags=-2.7327843e-009 walpha0=8.0653667e-012 wbeta0=1.2157547e-007 wint=1e-008 wk2=-7.9923454e-009 wketa=-7.1103921e-010 wkt1=-7.8619588e-009 wkt2=1.8375e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.3733463e-009 wr=1 wtvoff=0 wu0=7.2111957e-010 wua=6.5067587e-018 wub1=2.4014016e-026 wub=-1.7352055e-026 wuc=-9.5351961e-018 wute=1.8375e-008 wvoff=2.231366e-009 wvth0=-1.0403021e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.3 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.274905 alpha0=6.60855e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.88825 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=0.0059457 k3=0 k3b=0 keta=-0.02274975 kt1=-0.331385 kt1l=0 kt2=-0.021125 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.185545 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.03219475 ua1=1.675e-009 ua=-7.96735e-010 ub1=-2.5955e-018 ub=2.72215e-018 uc1=-5.6e-011 uc=9.86815e-011 ute=-1.3875 vbm=-3 version=4.5 vfbcv=-1 voff=-0.1251825 voffcv=0.005 voffl=0 vsat=92500 vth0=0.5916975 w0=5e-007 wags=2.05065e-009 walpha0=7.108185e-012 wbeta0=8.85675e-008 wint=1e-008 wk2=-7.716177e-009 wketa=-1.0021725e-009 wkt1=-6.32835e-009 wkt2=1.8375e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=7.37205e-009 wr=1 wtvoff=0 wu0=8.742825e-010 wua=8.59215e-018 wub1=3.7044e-026 wub=-2.91795e-026 wuc=-9.386685e-018 wute=1.8375e-008 wvoff=2.216025e-009 wvth0=-1.0793475e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.4 nmos a0=0.10668786 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.3531832 alpha0=2.618997e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=20.979752 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0039772727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.94866818 k2=0.037416157 k3=0 k3b=0 keta=-0.12161181 kt1=-0.37582777 kt1l=0 kt2=-0.014896384 ku0=0 kvsat=0 kvth0=0 la0=-1.5761839e-009 lags=-1.0591044e-008 lalpha0=-2.5821257e-013 lbeta0=-8.3833352e-008 ldelta=2.9210227e-009 level=54 lint=0 lk1=-9.1790218e-008 lk2=-3.4832437e-008 lketa=2.774773e-008 lkt1=1.529097e-008 lkt2=-3.0815037e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-7.3917648e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=3.7009358e-009 lua=3.665866e-016 lub1=2.2901987e-025 lub=-7.8888061e-026 luc=-3.141186e-017 lvoff=-8.5346442e-009 lvsat=0.0039725909 lvth0=-3.8570937e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=9.9275047e-016 pags=-1.3056615e-014 palpha0=-2.3504827e-020 paramchk=1 pbeta0=9.9761689e-014 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.45094152 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=3.3826512e-015 pketa=1.5971603e-015 pkt1=3.3480996e-015 pkt2=1.7961971e-015 ppclm=2.2974387e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.3091682e-016 pua=3.6449515e-024 pub1=-3.6790164e-032 pub=-2.3015752e-031 puc=-7.1059521e-024 pvag=0 pvoff=4.5598392e-015 pvsat=-1.9465696e-009 pvth0=1.8930389e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.033441305 ua1=1.675e-009 ua=-5.8760066e-010 ub1=-3.6336059e-018 ub=2.2723958e-018 uc1=-5.6e-011 uc=1.5510632e-010 ute=-1.435 vbm=-3 version=4.5 vfbcv=-1 voff=-0.080003796 voffcv=0.005 voffl=0 vsat=79409.091 vth0=0.6494457 w0=5e-007 wa0=-3.7462282e-009 wags=3.2518616e-008 walpha0=4.8463561e-014 wbeta0=-3.781252e-007 wint=1e-008 wk2=-1.2764722e-008 wketa=-3.293114e-009 wkt1=-6.9032982e-009 wkt2=-3.7034991e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.773173e-008 wr=1 wtvoff=0 wu0=8.8373727e-011 wua=1.9523816e-017 wub1=7.5856009e-026 wub=9.2037981e-026 wuc=-8.4901632e-019 wute=4.165e-008 wvoff=-1.720694e-008 wvsat=0.0098445454 wvth0=-2.2012593e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.5 nmos a0=0.9644116 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.43863251 alpha0=6.7595967e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.025956 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0015357143 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.76840415 k2=0.0076001761 k3=0 k3b=0 keta=-0.044144964 kt1=-0.40772797 kt1l=0 kt2=-0.031195536 ku0=0 kvsat=0 kvth0=0 la0=-4.175722e-007 lags=-5.2033959e-008 lalpha0=-2.2664034e-012 lbeta0=-1.0624202e-007 ldelta=4.1051786e-009 level=54 lint=0 lk1=-4.3621628e-009 lk2=-2.0371686e-008 lketa=-9.8236923e-009 lkt1=3.0762566e-008 lkt2=4.8235848e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=3.8780801e-008 lpdiblc2=8.6783475e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.7382792e-009 lua=6.3534043e-016 lub1=-1.6787717e-025 lub=-3.412717e-025 luc1=3.0374545e-017 luc=4.0251276e-018 lvoff=1.1009268e-008 lvsat=-0.004023075 lvth0=-1.6914157e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.3952024e-015 pags=-2.7575765e-014 palpha0=6.5383015e-020 paramchk=1 pbeta0=-2.8587971e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21857359 pdiblc1=0.39 pdiblc2=0.00138165 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=5.1909737e-015 pk2=-4.9643217e-015 pkt1=-1.5073657e-014 pkt2=-2.5647103e-015 ppclm=2.4333971e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.5085237e-016 pua=2.2200133e-023 pub1=-2.9340286e-032 pub=-2.3130267e-031 puc1=-1.4883527e-023 puc=-9.1474668e-024 pvag=0 pvoff=-6.4083562e-015 pvsat=4.7874593e-009 pvth0=-3.2623115e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.031302452 ua1=1.675e-009 ua=-1.1417323e-009 ub1=-2.8152615e-018 ub=2.813393e-018 uc1=-1.1862793e-010 uc=8.2040368e-011 ute=-1.435 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12030052 voffcv=0.005 voffl=0 vsat=95895 vth0=0.60479255 w0=5e-007 wa0=1.177386e-009 wags=6.2455008e-008 walpha0=-1.3481034e-013 wbeta0=4.170117e-007 wint=1e-008 wk1=-1.0703038e-008 wk2=4.4455318e-009 wkt1=3.1079706e-008 wkt2=5.2880625e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-2.0534997e-008 wr=1 wtvoff=0 wu0=1.2947795e-010 wua=-1.8734289e-017 wub1=6.0495435e-026 wub=9.439913e-026 wuc1=3.0687684e-017 wuc=3.3602922e-018 wute=4.165e-008 wvoff=5.4078955e-009 wvsat=-0.00404005 wvth0=-1.1383005e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.6 nmos a0=1.2324275 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.28413926 alpha0=9.079175e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.031764 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027306818 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79412996 k2=-0.0056941447 k3=0 k3b=0 keta=-0.021073023 kt1=-0.33925459 kt1l=0 kt2=-0.021820469 ku0=0 kvsat=0 kvth0=0 la0=-7.351711e-007 lags=1.3104055e-007 lalpha0=-1.018445e-010 lbeta0=-3.6681242e-006 ldelta=2.689142e-009 level=54 lint=0 lk1=-3.4847247e-008 lk2=-4.6179157e-009 lketa=-3.7163943e-008 lkt1=-5.0378387e-008 lkt2=-6.2858695e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=2.8319355e-008 lpdiblc2=1.7439086e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.433985e-009 lua=2.1582113e-016 lub1=7.0841414e-025 lub=-6.3545771e-025 luc1=-4.9742943e-017 luc=-1.4517602e-017 lute=3.4286561e-007 lvoff=1.297511e-008 lvth0=1.3266882e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=6.4659197e-014 palpha0=-1.0707464e-019 paramchk=1 pbeta0=-3.0240747e-014 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.22740181 pdiblc1=0.39 pdiblc2=0.00064234716 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-8.5010099e-015 pk2=2.7459718e-015 pkt1=2.468541e-014 pkt2=3.0800761e-015 ppclm=1.9533282e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.3496333e-015 pua=8.6354133e-024 pub1=-5.870065e-031 pub=8.5458111e-032 puc1=2.4374042e-023 puc=5.1476471e-024 pute=-1.6800415e-013 pvag=0 pvth0=-1.1771491e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.036511114 ua1=1.675e-009 ua=-7.8770753e-010 ub1=-3.5547478e-018 ub=3.0616512e-018 uc1=-5.1018233e-011 uc=9.7688241e-011 ute=-1.7243381 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12195946 voffcv=0.005 voffl=0 vsat=92500 vth0=0.57932332 w0=5e-007 wags=-1.5380403e-008 walpha0=1.072355e-014 wbeta0=2.0128262e-007 wint=1e-008 wk1=8.5137806e-010 wk2=-2.061045e-009 wkt1=-2.4722493e-009 wkt2=5.2452969e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.6483783e-008 wr=1 wtvoff=0 wu0=-1.3055311e-009 wua=-7.2872686e-018 wub1=5.3109983e-025 wub=-1.7290955e-025 wuc1=-2.4410658e-018 wuc=-8.703095e-018 wute=1.8342565e-007 wvth0=-4.2022626e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.7 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.297263 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.6644 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=-0.00615663 k3=0 k3b=0 keta=-0.024795 kt1=-0.3443 kt1l=0 kt2=-0.02245 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.230238 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.0363675 ua1=1.675e-009 ua=-7.66093e-010 ub1=-3.4838e-018 ub=2.99801e-018 uc1=-5.6e-011 uc=9.62343e-011 ute=-1.69 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.005 voffl=0 vsat=92500 vth0=0.580652 w0=5e-007 wags=-8.90477e-009 wbeta0=1.98254e-007 wint=1e-008 wk2=-1.7860353e-009 wkt2=8.33e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.452752e-008 wr=1 wtvoff=0 wu0=-1.170365e-009 wua=-6.42243e-018 wub1=4.72311e-025 wub=-1.643509e-025 wuc=-8.187557e-018 wute=1.666e-007 wvth0=-5.38118e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.8 nmos a0=0.10353977 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.27394573 alpha0=2.567968e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.141066 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0039772727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.94035419 k2=0.010689994 k3=0 k3b=0 keta=-0.12103166 kt1=-0.28213548 kt1l=0 kt2=-0.025353566 ku0=0 kvsat=0 kvth0=0 la0=-7.4193977e-010 lags=3.0120571e-008 lalpha0=-2.3346347e-013 ldelta=2.9210227e-009 level=54 lint=0 lk1=-8.7757932e-008 lk2=-2.7750003e-008 lketa=2.7466355e-008 lkt1=-9.299129e-009 lkt2=8.8905907e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.1937689e-006 lpclm=-8.9497813e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.5325411e-010 lua=2.3358646e-016 lub1=4.4342327e-025 lub=-3.051927e-025 luc1=4.5702115e-017 luc=-6.2506115e-017 lvoff=6.3595312e-010 lvoffcv=-1.0279677e-007 lvsat=-0.00031600155 lvth0=-5.1192629e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.46137913 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=-6.1503437e-014 palpha0=-5.2956251e-020 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.20348625 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-4.7984203e-015 pk2=-5.0454443e-015 pketa=1.9319955e-015 pkt1=3.2610317e-014 pkt2=-2.9287727e-015 pnoff=-1.420585e-012 ppclm=-5.4337375e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=3.8908244e-015 pua=1.6191512e-022 pub1=-2.9193021e-031 pub=3.9145008e-032 puc1=-5.4385517e-023 puc=2.9896211e-023 pvag=0 pvoff=-6.3531717e-015 pvoffcv=1.2232815e-013 pvsat=3.1568555e-009 pvth0=1.6912853e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.046929878 ua1=1.675e-009 ua=-6.3486383e-010 ub1=-5.3288522e-018 ub=3.762013e-018 uc1=-2.2422528e-010 uc=2.8720922e-010 ute=-1.5702841 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12420249 voffcv=0.21695209 voffl=0 vsat=93151.55 vth0=0.67826787 w0=5e-007 wags=1.2681121e-007 walpha0=1.0918815e-013 wbeta0=-5.7008843e-007 wint=1e-008 wk1=9.8936502e-009 wk2=1.9039412e-008 wketa=-3.983496e-009 wkt1=-1.1839713e-007 wkt2=8.7405474e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=2.9290412e-006 wpclm=2.7674005e-007 wr=1 wtvoff=0 wu0=-1.5963029e-008 wua=7.5766988e-017 wub1=2.0931991e-024 wub=-1.6806064e-024 wuc1=2.0018808e-016 wuc=-1.5805146e-016 wute=2.0263807e-007 wvoff=3.538951e-008 wvoffcv=-2.5222299e-007 wvsat=-0.0065089804 wvth0=-5.631097e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.9 nmos a0=0.57333915 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.62982962 alpha0=6.6463107e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.044461 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0015357143 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.016364333 k3=0 k3b=0 keta=-0.044144964 kt1=-0.30287445 kt1l=0 kt2=-0.021815574 ku0=0 kvsat=0 kvth0=0 la0=-2.2859464e-007 lags=-1.4248312e-007 lalpha0=-2.2114597e-012 lbeta0=4.6853149e-008 ldelta=4.1051786e-009 level=54 lint=0 lk2=-3.0502058e-008 lketa=-9.8236923e-009 lkt1=7.5927144e-010 lkt2=-8.2686693e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=6.5837837e-008 lpdiblc2=8.6783475e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.2020412e-009 lua=3.7138544e-016 lub1=-6.6136013e-025 lub=-1.6300526e-025 luc1=7.2679686e-018 luc=4.9517784e-019 lvoff=-9.7549306e-009 lvth0=-9.5240796e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.262785e-013 pags=8.0058731e-014 paramchk=1 pbeta0=-4.6806296e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.049284973 pdiblc1=0.39 pdiblc2=0.00138165 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=7.0908211e-015 pkt1=2.0630263e-014 pkt2=4.1593273e-015 ppclm=-7.8639014e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=2.8727087e-016 pua=3.3630657e-022 pub1=5.5790443e-031 pub=-4.4343974e-031 puc1=1.2613299e-023 puc=-4.9468266e-024 pvag=0 pvoff=1.830104e-014 pvth0=-1.2056503e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.038581863 ua1=1.675e-009 ua=-9.1898543e-010 ub1=-3.0509483e-018 ub=3.468843e-018 uc1=-1.4497962e-010 uc=1.5730964e-010 ute=-1.5702841 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10277799 voffcv=0.005 voffl=0 vsat=92500 vth0=0.59235333 w0=5e-007 wa0=4.665536e-007 wags=-1.6506955e-007 wbeta0=3.9498984e-007 wint=1e-008 wk2=-5.9838153e-009 wkt1=-9.3695983e-008 wkt2=-5.8740916e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.8091845e-007 wr=1 wtvoff=0 wu0=-8.5330215e-009 wua=-2.8380301e-016 wub1=3.4096267e-025 wub=-6.8558634e-025 wuc1=6.2046194e-017 wuc=-8.6210147e-017 wute=2.0263807e-007 wvoff=-1.5443916e-008 wvth0=3.4196621e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.10 nmos a0=1.1740916 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26765145 alpha0=9.0800762e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.507475 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027306818 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79742159 k2=-0.0074261153 k3=0 k3b=0 keta=-0.021073023 kt1=-0.31501857 kt1l=0 kt2=-0.016816848 ku0=0 kvsat=0 kvth0=0 la0=-9.4048631e-007 lags=2.8669802e-007 lalpha0=-1.0193448e-010 lbeta0=-4.0568183e-006 ldelta=2.689142e-009 level=54 lint=0 lk1=-4.504374e-008 lk2=-2.3103764e-009 lketa=-3.7163943e-008 lkt1=1.5150046e-008 lkt2=-6.7503577e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.5263937e-007 lpclm=-1.5218617e-007 lpdiblc2=1.7439086e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.9271691e-009 lua1=2.5643414e-017 lua=2.4275299e-016 lub1=-1.7294942e-024 lub=1.6734577e-025 luc1=-1.1139275e-016 luc=6.3166633e-017 lute=-2.7273401e-008 lvoff=1.297511e-008 lvoffcv=8.3951653e-008 lvth0=7.2824411e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1288096 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.4432511e-013 pags=-1.205732e-013 paramchk=1 pbeta0=4.3230522e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23327148 pdiblc1=0.39 pdiblc2=0.00064234716 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=3.632817e-015 pkt1=-5.3293425e-014 pkt2=3.632817e-015 pnoff=1.8164085e-013 ppclm=2.3433486e-013 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-2.65014e-015 pua1=-3.0515663e-023 pua=-2.3413506e-023 pub1=2.3141044e-030 pub=-8.6987803e-031 puc1=9.7737308e-023 puc=-8.7296592e-023 pute=2.7246128e-013 pvag=0 pvoffcv=-9.9902467e-014 pvth0=-4.6500058e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040501587 ua1=1.65336e-009 ua=-8.1043485e-010 ub1=-2.1495693e-018 ub=3.1900657e-018 uc1=-4.4843991e-011 uc=1.0442234e-010 ute=-1.5472686 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12195946 voffcv=-0.065845277 voffl=0 vsat=92500 vth0=0.57817062 w0=5e-007 wa0=6.9419757e-008 wags=4.2400941e-009 wbeta0=-3.6481453e-007 wint=1e-008 wk1=-3.0656684e-009 wkt1=-3.1313123e-008 wkt2=-5.4297792e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.5328342e-007 wpclm=-2.3468689e-008 wr=1 wtvoff=0 wu0=-6.0541938e-009 wua1=2.5751614e-017 wua=1.9758233e-017 wub1=-1.1410626e-024 wub=-3.2572281e-025 wuc1=-9.7884135e-018 wuc=-1.6716674e-017 wute=-2.7287058e-008 wvoffcv=8.430588e-008 wvth0=-2.8305468e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.11 nmos a0=1.0799017 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29636432 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.101184 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79291046 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31350128 kt1l=0 kt2=-0.017492898 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1135227 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040694593 ua1=1.6559282e-009 ua=-7.8612308e-010 ub1=-2.3227785e-018 ub=3.2068255e-018 uc1=-5.6e-011 uc=1.1074849e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.0574375 voffl=0 vsat=92500 vth0=0.57889996 w0=5e-007 wa0=9.3888972e-008 wags=-7.8353386e-009 wbeta0=-3.2151907e-007 wint=1e-008 wk1=-2.7018409e-009 wkt1=-3.6650472e-008 wkt2=-5.0659517e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.3509204e-007 wr=1 wtvoff=0 wu0=-6.3196059e-009 wua1=2.2695464e-017 wua=1.7413365e-017 wub1=-9.0930456e-025 wub=-4.1284129e-025 wuc=-2.5459447e-017 wvoffcv=7.4300625e-008 wvth0=-3.2962459e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.12 nmos a0=0.13050819 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.45484419 alpha0=2.5788977e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=2.07e-010 cgidl=0.5 cgsl=9e-011 cgso=2.07e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0039772727 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.94134454 k2=0.012595841 k3=0 k3b=0 keta=-0.11802055 kt1=-0.29398705 kt1l=0 kt2=-0.024478636 ku0=0 kvsat=0 kvth0=0 la0=-1.3821621e-008 lags=-5.7615181e-008 lalpha0=-2.387644e-013 ldelta=2.9210227e-009 level=54 lint=0 lk1=-8.8238255e-008 lk2=-2.8255053e-008 lketa=2.6005966e-008 lkt1=-6.034833e-009 lkt2=5.9588864e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.0515682e-006 lpclm=-1.4388958e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=5.4272602e-010 lua=2.4979418e-016 lub1=4.1420102e-025 lub=-3.0127428e-025 luc1=4.0258119e-017 luc=-5.9513501e-017 lvoffcv=-9.0551705e-008 lvth0=-4.9499651e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.16818182 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.3066601e-013 pags=8.1497672e-013 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23118796 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pketa=1.6521288e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.045331977 ua1=1.675e-009 ua=-6.2727955e-010 ub1=-5.1193227e-018 ub=3.5937841e-018 uc1=-2.0418643e-010 uc=2.7138825e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.19170454 voffl=0 vsat=92500 vth0=0.67263114 w0=5e-007 wa0=-2.6941446e-007 wags=-1.6803644e-006 wint=1e-008 wketa=-3.4064511e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.13 nmos a0=0.62004121 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.61330614 alpha0=6.6463107e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0015357143 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.015765353 k3=0 k3b=0 keta=-0.044144964 kt1=-0.31225343 kt1l=0 kt2=-0.022403571 ku0=0 kvsat=0 kvth0=0 la0=-2.5124514e-007 lags=-1.3446923e-007 lalpha0=-2.2114597e-012 ldelta=4.1051786e-009 level=54 lint=0 lk2=-2.9792266e-008 lketa=-9.8236923e-009 lkt1=2.8243629e-009 lkt2=-4.1051786e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=6.505066e-008 lpdiblc2=8.6783475e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.230797e-009 lua=4.0504976e-016 lub1=-6.0551384e-025 lub=-2.0739362e-025 luc1=8.5305611e-018 lvoff=-7.9229946e-009 lvth0=-1.0730937e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.067394929 pdiblc1=0.39 pdiblc2=0.00138165 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.037727707 ua1=1.675e-009 ua=-9.4739414e-010 ub1=-3.0168179e-018 ub=3.4002157e-018 uc1=-1.3876879e-010 uc=1.4868e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10432393 voffcv=0.005 voffl=0 vsat=92500 vth0=0.59269564 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.14 nmos a0=1.1810406 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26807588 alpha0=9.0800762e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.470957 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=7.7e-011 cgidl=0.5 cgsl=9e-011 cgso=7.7e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027306818 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79711472 k2=-0.0074261153 k3=0 k3b=0 keta=-0.021073023 kt1=-0.31815301 kt1l=0 kt2=-0.017360369 ku0=0 kvsat=0 kvth0=0 la0=-9.1602935e-007 lags=2.7462863e-007 lalpha0=-1.0193448e-010 lbeta0=-4.0135445e-006 ldelta=2.689142e-009 level=54 lint=0 lk1=-4.4680095e-008 lk2=-2.3103764e-009 lketa=-3.7163943e-008 lkt1=9.8153685e-009 lkt2=-6.3867124e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.344571e-007 lpclm=-1.2872923e-007 lpdiblc2=1.7439086e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.6618898e-009 lua1=2.2588793e-017 lua=2.404093e-016 lub1=-1.4978521e-024 lub=8.027089e-026 luc1=-1.0160923e-016 luc=5.4428235e-017 lvoff=1.297511e-008 lvoffcv=7.3951406e-008 lvth0=6.8169751e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1134659 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23092226 pdiblc1=0.39 pdiblc2=0.00064234716 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.039895561 ua1=1.6559377e-009 ua=-8.0845705e-010 ub1=-2.2637898e-018 ub=3.1574609e-018 uc1=-4.5823812e-011 uc=1.02749e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12195946 voffcv=-0.05740625 voffl=0 vsat=92500 vth0=0.57788728 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.model nmos_3p3.15 nmos a0=1.0893 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29558 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.069 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9e-011 cgdo=2.07e-010 cgidl=0.5 cgsl=9e-011 cgso=2.07e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79264 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31717 kt1l=0 kt2=-0.018 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.6e-009 toxm=8e-009 toxp=7.6e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040062 ua1=1.6582e-009 ua=-7.8438e-010 ub1=-2.4138e-018 ub=3.1655e-018 uc1=-5.6e-011 uc=1.082e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.05 voffl=0 vsat=92500 vth0=0.57857 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.5e-008 xpart=0 xtis=3 xw=1e-008
.subckt nplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 r_rsh0='rsh_nplus_u_m' r_dw=-5e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.36e-3 r_tc2=6.5e-7 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model np_junction d cj=0.00096797 level=2
d1 3 1 np_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends nplus_u_m1
.endl nmos_3p3_f

.lib nmos_3p3_s
.subckt nmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.007148
.param par_k=0.007008
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b nplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b nplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b nmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model nmos_3p3.0 nmos a0=0.11164211 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.33078713 alpha0=2.689932e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=19.906217 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0032954546 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.97009364 k2=0.057112207 k3=0 k3b=0 keta=-0.15224321 kt1=-0.46042018 kt1l=0 kt2=-0.024751234 ku0=0 kvsat=0 kvth0=0 la0=-3.216124e-009 lags=-1.7784597e-008 lalpha0=-3.3259243e-013 lbeta0=1.3969208e-007 ldelta=3.4528409e-009 level=54 lint=0 lk1=-1.0850207e-007 lk2=-4.4586066e-008 lketa=4.1863427e-008 lkt1=4.4736487e-008 lkt2=1.327864e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-5.0349819e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.9752231e-009 lua=7.4602352e-016 lub1=3.0544077e-025 lub=-8.4745491e-025 luc1=-3.9362386e-018 luc=-6.5971448e-017 lute=9.3719968e-008 lvoff=4.1027149e-009 lvsat=-0.002811599 lvth0=-4.1963855e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.7614949e-015 pags=-1.2329143e-014 palpha0=-1.3787144e-020 paramchk=1 pbeta0=8.809677e-016 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.38126164 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=5.4388743e-015 pketa=-2.4490902e-015 pkt1=-8.7347947e-015 pkt2=-2.9952902e-016 ppclm=8.6466979e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-6.5742214e-016 pua=-1.428335e-022 pub1=-5.8033747e-032 pub=9.3519126e-032 puc1=1.8500322e-024 puc=5.4982075e-024 pute=-4.4048385e-014 pvag=0 pvoff=-1.4998475e-015 pvsat=1.3214515e-009 pvth0=4.4048385e-016 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.02365998 ua1=1.675e-009 ua=-1.2009004e-009 ub1=-4.1897925e-018 ub=3.4181442e-018 uc1=-4.2656818e-011 uc=2.2972174e-010 ute=-1.5659091 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12611751 voffcv=0.005 voffl=0 vsat=82709.416 vth0=0.78102964 w0=5e-007 wa0=-5.9711692e-009 wags=4.5802637e-008 walpha0=4.6736083e-014 wbeta0=1.2873117e-007 wint=1e-008 wk2=-1.8436862e-008 wketa=7.8363649e-009 wkt1=3.0709777e-008 wkt2=1.0153526e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=1.8707045e-008 wr=1 wtvoff=0 wu0=4.3500625e-009 wua=2.6594489e-016 wub1=3.1727957e-025 wub=-3.9003587e-025 wuc1=-6.2712955e-018 wuc=-3.0846577e-017 wute=1.0147727e-007 wvoff=5.0842288e-009 wvsat=-0.00033342533 wvth0=-1.335093e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.1 nmos a0=1.0928896 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.48554907 alpha0=6.6270642e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=22.618932 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0013214286 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.74623593 k2=0.024093133 k3=0 k3b=0 keta=-0.028668661 kt1=-0.33899638 kt1l=0 kt2=-0.020292087 ku0=0 kvsat=0 kvth0=0 la0=-5.0855857e-007 lags=-9.7486997e-008 lalpha0=-2.3602156e-012 lbeta0=-1.2573561e-006 ldelta=4.4694643e-009 level=54 lint=0 lk1=6.7846468e-009 lk2=-2.7581243e-008 lketa=-2.1777465e-008 lkt1=-1.7796768e-008 lkt2=-9.6859676e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=1.0221633e-007 lpdiblc2=9.4484475e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.8540296e-009 lua=8.0247348e-016 lub1=-4.1622844e-025 lub=-6.8218008e-025 luc1=5.0951893e-018 luc=8.7468885e-018 lvoff=-2.9137715e-009 lvsat=0.0020112589 lvth0=-2.4499049e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.3890942e-014 pags=-9.6046138e-015 palpha0=1.7846507e-020 paramchk=1 pbeta0=2.3804846e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.085016691 pdiblc1=0.39 pdiblc2=0.00133635 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=-2.6453883e-015 pketa=5.2085573e-015 pkt1=8.3644811e-015 pkt2=2.4517566e-016 ppclm=-2.7853095e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.1868212e-015 pua=-2.8870859e-023 pub1=7.9083403e-032 pub=-9.5555786e-032 puc1=-2.394739e-024 puc=-1.160405e-023 pvag=0 pvoff=3.1074589e-016 pvsat=1.9956158e-009 pvth0=-5.4736891e-016 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.02972055 ua1=1.675e-009 ua=-1.310512e-009 ub1=-2.788493e-018 ub=3.0972222e-018 uc1=-6.0193571e-011 uc=8.4637593e-011 ute=-1.3839286 vbm=-3 version=4.5 vfbcv=-1 voff=-0.11249326 voffcv=0.005 voffl=0 vsat=73344.643 vth0=0.7471174 w0=5e-007 wa0=-4.894097e-008 wags=4.0512289e-008 walpha0=-1.4688483e-014 wbeta0=-3.3178823e-007 wint=1e-008 wk2=-2.7392647e-009 wketa=-7.0328534e-009 wkt1=-2.4927001e-009 wkt2=-4.2326378e-011 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=4.0905118e-008 wr=1 wtvoff=0 wu0=7.6900741e-010 wua=4.4658224e-017 wub1=5.1032672e-026 wub=-2.2900119e-026 wuc1=1.9709786e-018 wuc=2.3616893e-018 wute=1.5946429e-008 wvoff=1.5685135e-009 wvsat=-0.0016424821 wvth0=-1.1432769e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.2 nmos a0=1.2256909 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.25735343 alpha0=7.6135347e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.225975 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027238636 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79599981 k2=0.0048675395 k3=0 k3b=0 keta=-0.019679504 kt1=-0.32971157 kt1l=0 kt2=-0.021089286 ku0=0 kvsat=0 kvth0=0 la0=-6.6991215e-007 lags=1.7977071e-007 lalpha0=-8.6812779e-011 lbeta0=-3.2099126e-006 ldelta=2.7655057e-009 level=54 lint=0 lk1=-5.3678465e-008 lk2=-4.2221469e-009 lketa=-3.269929e-008 lkt1=-2.9077811e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=-2.465794e-008 lpdiblc2=1.7934304e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.5461646e-009 lua=2.0053373e-016 lub1=-7.505138e-025 lub=-2.4989307e-025 luc=-6.9419625e-018 lvoff=1.3634437e-008 lvth0=-3.6588628e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-4.0483744e-014 pags=4.2627001e-014 palpha0=-8.5298102e-018 paramchk=1 pbeta0=-2.9414659e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.18943996 pdiblc1=0.39 pdiblc2=0.00063792557 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=2.4610412e-015 pketa=-2.5943994e-015 pkt1=1.3666571e-014 ppclm=4.4545348e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.3648931e-015 pua=1.8583714e-023 pub1=1.1611514e-031 pub=-1.0539885e-031 puc=1.3234392e-024 pvag=0 pvoff=-1.3670981e-016 pvth0=-3.4794852e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032519064 ua1=1.675e-009 ua=-8.1508834e-010 ub1=-2.513361e-018 ub=2.7414305e-018 uc1=-5.6e-011 uc=9.7550228e-011 ute=-1.3839286 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12611319 voffcv=0.005 voffl=0 vsat=75000 vth0=0.72996498 w0=5e-007 wa0=4.0423109e-009 wags=-2.4766942e-009 walpha0=7.0204199e-012 wbeta0=1.0623239e-007 wint=1e-008 wk2=-6.9420874e-009 wketa=-6.1066685e-010 wkt1=-6.8565602e-009 wkt2=1.5946429e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=1.9498441e-009 wr=1 wtvoff=0 wu0=6.2244619e-010 wua=5.600962e-018 wub1=2.0553877e-026 wub=-1.4798829e-026 wuc=-8.2782193e-018 wute=1.5946429e-008 wvoff=1.9367898e-009 wvth0=-9.0195048e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.3 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.27530357 alpha0=6.7467071e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.905464 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=0.0044459571 k3=0 k3b=0 keta=-0.022944536 kt1=-0.332615 kt1l=0 kt2=-0.021089286 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.18697786 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032364679 ua1=1.675e-009 ua=-7.95065e-010 ub1=-2.5883e-018 ub=2.7164786e-018 uc1=-5.6e-011 uc=9.6857071e-011 ute=-1.3839286 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12475179 voffcv=0.005 voffl=0 vsat=75000 vth0=0.72959964 w0=5e-007 wags=1.7796214e-009 walpha0=6.1687164e-012 wbeta0=7.6861786e-008 wint=1e-008 wk2=-6.6963519e-009 wketa=-8.6971821e-010 wkt1=-5.49195e-009 wkt2=1.5946429e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=6.3977071e-009 wr=1 wtvoff=0 wu0=7.5873107e-010 wua=7.45655e-018 wub1=3.2148e-026 wub=-2.5322929e-026 wuc=-8.1460736e-018 wute=1.5946429e-008 wvoff=1.9231393e-009 wvth0=-9.3669321e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.4 nmos a0=0.10691933 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.35687524 alpha0=2.6811189e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=20.985552 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0032954546 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.97009364 k2=0.045081757 k3=0 k3b=0 keta=-0.12821436 kt1=-0.37966054 kt1l=0 kt2=-0.014318515 ku0=0 kvsat=0 kvth0=0 la0=-1.8229027e-009 lags=-1.304868e-008 lalpha0=-3.0617722e-013 lbeta0=-9.5051778e-008 ldelta=3.4528409e-009 level=54 lint=0 lk1=-1.0850207e-007 lk2=-4.1037083e-008 lketa=3.2864396e-008 lkt1=1.8210678e-008 lkt2=-3.5697146e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-8.6444043e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.3613327e-009 lua=4.3347724e-016 lub1=2.6922491e-025 lub=-1.0258242e-025 luc=-3.7418989e-017 lvoff=-9.9036356e-009 lvsat=0.0046169416 lvth0=-4.5516631e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.1066809e-015 pags=-1.4555024e-014 palpha0=-2.6202298e-020 paramchk=1 pbeta0=1.1121058e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.46740308 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=3.7708524e-015 pketa=1.7804543e-015 pkt1=3.7323356e-015 pkt2=2.0023329e-015 ppclm=2.5610983e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.6889363e-016 pua=4.0632548e-024 pub1=-4.1012292e-032 pub=-2.5657094e-031 puc=-7.9214482e-024 pvag=0 pvoff=5.0831372e-015 pvsat=-2.1699625e-009 pvth0=2.1102886e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032583121 ua1=1.675e-009 ua=-6.7252796e-010 ub1=-3.6841668e-018 ub=2.2958092e-018 uc1=-5.6e-011 uc=1.6246617e-010 ute=-1.4335714 vbm=-3 version=4.5 vfbcv=-1 voff=-0.078638354 voffcv=0.005 voffl=0 vsat=61335.065 vth0=0.79767867 w0=5e-007 wa0=-3.7514606e-009 wags=3.3541222e-008 walpha0=5.0878248e-014 wbeta0=-3.7855616e-007 wint=1e-008 wk2=-1.2782551e-008 wketa=-3.4571927e-009 wkt1=-7.2472535e-009 wkt2=-3.8880251e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-2.1779432e-008 wr=1 wtvoff=0 wu0=1.5618588e-010 wua=1.7609833e-017 wub1=7.9635518e-026 wub=1.3746161e-025 wuc=7.6353972e-019 wute=3.9278571e-008 wvoff=-1.7230974e-008 wvsat=0.0097125195 wvth0=-2.1175971e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.5 nmos a0=0.98625128 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.44354017 alpha0=6.8731595e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.046316 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0013214286 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.76825545 k2=0.0088249226 k3=0 k3b=0 keta=-0.043632179 kt1=-0.40824074 kt1l=0 kt2=-0.031261352 ku0=0 kvsat=0 kvth0=0 la0=-4.5467886e-007 lags=-5.7681118e-008 lalpha0=-2.4650781e-012 lbeta0=-1.2634537e-007 ldelta=4.4694643e-009 level=54 lint=0 lk1=-4.5554057e-009 lk2=-2.2364814e-008 lketa=-1.0695428e-008 lkt1=3.292948e-008 lkt2=5.1558463e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=4.3130841e-008 lpdiblc2=9.4484475e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=5.1456432e-009 lua=6.9254834e-016 lub1=-1.8386993e-025 lub=-3.8019306e-025 luc1=3.2514127e-017 luc=4.040715e-018 lvoff=1.1746901e-008 lvsat=-0.0042012964 lvth0=-1.8536912e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.432522e-015 pags=-2.8313377e-014 palpha0=6.7131915e-020 paramchk=1 pbeta0=-2.9352658e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21580136 pdiblc1=0.39 pdiblc2=0.00133635 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=5.3298247e-015 pk2=-5.0971101e-015 pkt1=-1.5476856e-014 pkt2=-2.6333126e-015 ppclm=2.498487e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.6023716e-016 pua=2.2793954e-023 pub1=-3.0125096e-032 pub=-2.3748968e-031 puc1=-1.528164e-023 puc=-9.3921482e-024 pvag=0 pvoff=-6.5797704e-015 pvsat=4.9155168e-009 pvth0=-3.3495736e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.031060188 ua1=1.675e-009 ua=-1.1755786e-009 ub1=-2.804371e-018 ub=2.834859e-018 uc1=-1.1913423e-010 uc=8.1961894e-011 ute=-1.4335714 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12067823 voffcv=0.005 voffl=0 vsat=78457.857 vth0=0.74529086 w0=5e-007 wa0=1.1790305e-009 wags=6.0256471e-008 walpha0=-1.3035323e-013 wbeta0=4.0734123e-007 wint=1e-008 wk1=-1.0349174e-008 wk2=4.4367941e-009 wkt1=3.0052147e-008 wkt2=5.1132283e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-2.0563679e-008 wr=1 wtvoff=0 wu0=1.393772e-010 wua=-1.8760456e-017 wub1=5.8495332e-026 wub=1.0041062e-025 wuc1=2.9673087e-017 wuc=3.6192678e-018 wute=3.9278571e-008 wvoff=5.4154489e-009 wvsat=-0.0040456929 wvth0=-1.0574296e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.6 nmos a0=1.2342915 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.28327385 alpha0=9.1050349e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.04797 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027238636 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79424825 k2=-0.0057533677 k3=0 k3b=0 keta=-0.020978796 kt1=-0.3392138 kt1l=0 kt2=-0.021786808 ku0=0 kvsat=0 kvth0=0 la0=-7.5604777e-007 lags=1.3704246e-007 lalpha0=-1.0474036e-010 lbeta0=-3.7733547e-006 ldelta=2.7655057e-009 level=54 lint=0 lk1=-3.6136665e-008 lk2=-4.6521909e-009 lketa=-3.8219289e-008 lkt1=-5.0938244e-008 lkt2=-6.3557247e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=2.9812546e-008 lpdiblc2=1.7934304e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.4270997e-009 lua=2.2225441e-016 lub1=7.0782525e-025 lub=-6.5048842e-025 luc1=-5.0295738e-017 luc=-1.4748284e-017 lute=3.4667589e-007 lvoff=1.3343565e-008 lvth0=1.3228401e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=6.2709277e-014 palpha0=-1.0384561e-019 paramchk=1 pbeta0=-2.932878e-014 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.22676292 pdiblc1=0.39 pdiblc2=0.00063792557 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-8.244646e-015 pk2=2.6631619e-015 pkt1=2.3940975e-014 pkt2=2.9871906e-015 ppclm=1.894422e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.3089326e-015 pua=8.3749962e-024 pub1=-5.6930421e-031 pub=8.2880961e-032 puc1=2.3638997e-023 puc=4.9924102e-024 pute=-1.6293767e-013 pvag=0 pvth0=-1.1416499e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.036469853 ua1=1.675e-009 ua=-7.8850544e-010 ub1=-3.5382765e-018 ub=3.0573243e-018 uc1=-5.0977959e-011 uc=9.7426091e-011 ute=-1.7189014 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12199236 voffcv=0.005 voffl=0 vsat=75000 vth0=0.71914657 w0=5e-007 wags=-1.4659294e-008 walpha0=1.0369007e-014 wbeta0=1.8989449e-007 wint=1e-008 wk1=8.2322976e-010 wk2=-1.950261e-009 wkt1=-2.3905117e-009 wkt2=4.8729978e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.559195e-008 wr=1 wtvoff=0 wu0=-1.2344251e-009 wua=-6.893001e-018 wub1=5.0226415e-025 wub=-1.6326892e-025 wuc1=-2.3603592e-018 wuc=-8.2198748e-018 wute=1.7338365e-007 wvth0=-3.9348514e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.7 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29695757 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.6712 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=-0.00621789 k3=0 k3b=0 keta=-0.024795 kt1=-0.3443 kt1l=0 kt2=-0.022421429 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.22973971 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.036327357 ua1=1.675e-009 ua=-7.6631329e-010 ub1=-3.4676e-018 ub=2.9923729e-018 uc1=-5.6e-011 uc=9.5953471e-011 ute=-1.6842857 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.005 voffl=0 vsat=75000 vth0=0.72046743 w0=5e-007 wags=-8.3977586e-009 wbeta0=1.86966e-007 wint=1e-008 wk2=-1.6843437e-009 wkt2=7.8557143e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.3700366e-008 wr=1 wtvoff=0 wu0=-1.1037279e-009 wua=-6.0567557e-018 wub1=4.45419e-025 wub=-1.5499324e-025 wuc=-7.7213816e-018 wute=1.5711429e-007 wvth0=-5.0747914e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.8 nmos a0=0.10371296 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26715255 alpha0=2.622667e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.140107 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0032954546 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.96085697 k2=0.017201346 k3=0 k3b=0 keta=-0.12745025 kt1=-0.28017689 kt1l=0 kt2=-0.025545233 ku0=0 kvsat=0 kvth0=0 la0=-8.7702159e-010 lags=3.5482186e-008 lalpha0=-2.7607448e-013 ldelta=3.4528409e-009 level=54 lint=0 lk1=-1.0374519e-007 lk2=-3.2812362e-008 lketa=3.247088e-008 lkt1=-1.0927331e-008 lkt2=1.045102e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.4082882e-006 lpclm=-1.0687288e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.8889394e-010 lua=2.7643655e-016 lub1=5.2357491e-025 lub=-3.6068e-025 luc1=5.3914751e-017 luc=-7.3826884e-017 lvoff=7.3910414e-010 lvoffcv=-1.2126927e-007 lvsat=-0.00036725671 lvth0=-6.047942e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.73454029 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=-7.1336137e-014 palpha0=-6.1422492e-020 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.2060622 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-5.5655552e-015 pk2=-5.8520714e-015 pketa=2.2408683e-015 pkt1=3.7823806e-014 pkt2=-3.3970025e-015 pnoff=-1.6476972e-012 ppclm=-6.302442e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=4.5128597e-015 pua=1.8780087e-022 pub1=-3.3860178e-031 pub=4.5403213e-032 puc1=-6.3080258e-023 puc=3.4675789e-023 pvag=0 pvoff=-7.3688683e-015 pvoffcv=1.4188504e-013 pvsat=3.6615494e-009 pvth0=1.9616751e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.046865722 ua1=1.675e-009 ua=-6.8932314e-010 ub1=-5.4287188e-018 ub=3.8304076e-018 uc1=-2.3453481e-010 uc=3.0152161e-010 ute=-1.5699432 vbm=-3 version=4.5 vfbcv=-1 voff=-0.1242889 voffcv=0.2404743 voffl=0 vsat=75713.12 vth0=0.83011576 w0=5e-007 wags=1.3851677e-007 walpha0=1.1926697e-013 wbeta0=-5.5938498e-007 wint=1e-008 wk1=1.0806903e-008 wk2=1.983753e-008 wketa=-4.3512005e-009 wkt1=-1.2364312e-007 wkt2=9.247235e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=3.1994121e-006 wpclm=2.839894e-007 wr=1 wtvoff=0 wu0=-1.6554457e-008 wua=3.7260197e-017 wub1=2.1207614e-024 wub=-1.6580185e-024 wuc1=2.0888573e-016 wuc=-1.6193132e-016 wute=1.9883352e-007 wvoff=3.618017e-008 wvoffcv=-2.7550493e-007 wvsat=-0.0071098048 wvth0=-5.9127366e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.9 nmos a0=0.58607632 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.63698234 alpha0=6.7617464e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.042721 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0013214286 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.017945817 k3=0 k3b=0 keta=-0.043632179 kt1=-0.30307353 kt1l=0 kt2=-0.02178266 ku0=0 kvsat=0 kvth0=0 la0=-2.4929415e-007 lags=-1.5498016e-007 lalpha0=-2.4077004e-012 lbeta0=5.0153484e-008 ldelta=4.4694643e-009 level=54 lint=0 lk2=-3.3195765e-008 lketa=-1.0695428e-008 lkt1=8.6443502e-010 lkt2=-8.9262312e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=7.1665757e-008 lpdiblc2=9.4484475e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.5754485e-009 lua=4.0495747e-016 lub1=-7.1902608e-025 lub=-1.7828226e-025 luc1=7.9360174e-018 luc=5.3005815e-019 lvoff=-1.0587044e-008 lvth0=-1.0391311e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.4173263e-013 pags=8.5526499e-014 paramchk=1 pbeta0=-5.0003024e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.046153372 pdiblc1=0.39 pdiblc2=0.00133635 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=7.5751026e-015 pkt1=2.2039247e-014 pkt2=4.4433966e-015 ppclm=-8.4009819e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=3.068906e-016 pua=3.5927528e-022 pub1=5.960076e-031 pub=-4.7372533e-031 puc1=1.3474748e-023 puc=-5.2846797e-024 pvag=0 pvoff=1.9550945e-014 pvth0=-1.2879926e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.038348141 ua1=1.675e-009 ua=-9.3887833e-010 ub1=-3.0159014e-018 ub=3.4762372e-018 uc1=-1.4525572e-010 uc=1.5713919e-010 ute=-1.5699432 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10229638 voffcv=0.005 voffl=0 vsat=75000 vth0=0.73285729 w0=5e-007 wa0=4.6938374e-007 wags=-1.6607087e-007 wbeta0=4.1154752e-007 wint=1e-008 wk2=-6.2346523e-009 wkt1=-9.2993492e-008 wkt2=-5.976841e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.7792447e-007 wr=1 wtvoff=0 wu0=-8.387527e-009 wua=-2.9569982e-016 wub1=3.0598585e-025 wub=-6.5000193e-025 wuc1=6.0235233e-017 wuc=-8.4338174e-017 wute=1.9883352e-007 wvoff=-1.6091313e-008 wvth0=3.9729778e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.10 nmos a0=1.1765919 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26693219 alpha0=9.1059211e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.517146 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027238636 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79753063 k2=-0.0074202574 k3=0 k3b=0 keta=-0.020978796 kt1=-0.31510943 kt1l=0 kt2=-0.016808883 ku0=0 kvsat=0 kvth0=0 la0=-9.6677061e-007 lags=2.9463078e-007 lalpha0=-1.0482912e-010 lbeta0=-4.1712719e-006 ldelta=2.7655057e-009 level=54 lint=0 lk1=-4.6316563e-008 lk2=-2.3759842e-009 lketa=-3.8219289e-008 lkt1=1.5488057e-008 lkt2=-6.9357625e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.5665961e-007 lpclm=-1.5610238e-007 lpdiblc2=1.7934304e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.9773099e-009 lua1=2.6318815e-017 lua=2.4960595e-016 lub1=-1.774603e-024 lub=1.7059289e-025 luc1=-1.1438687e-016 luc=6.4809343e-017 lute=-2.7576491e-008 lvoff=1.3343565e-008 lvoffcv=8.6162786e-008 lvth0=7.4811957e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.128938 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.4654573e-013 pags=-1.2166906e-013 paramchk=1 pbeta0=4.3623435e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23361686 pdiblc1=0.39 pdiblc2=0.00063792557 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=3.6658349e-015 pkt1=-5.3777798e-014 pkt2=3.6658349e-015 pnoff=1.8329175e-013 ppclm=2.3646468e-013 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-2.6742266e-015 pua1=-3.0793013e-023 pua=-2.3626306e-023 pub1=2.3351368e-030 pub=-8.7778417e-031 puc1=9.8625623e-023 puc=-8.8090013e-023 pute=2.7493762e-013 pvag=0 pvoffcv=-1.0081046e-013 pvth0=-4.6922687e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040486527 ua1=1.6533384e-009 ua=-8.1101699e-010 ub1=-2.1471138e-018 ub=3.1890972e-018 uc1=-4.4578445e-011 uc=1.0423443e-010 ute=-1.5472465 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12199236 voffcv=-0.065915874 voffl=0 vsat=75000 vth0=0.71814741 w0=5e-007 wa0=6.7508553e-008 wags=4.4604535e-009 wbeta0=-3.5904062e-007 wint=1e-008 wk1=-3.0171481e-009 wkt1=-3.0592631e-008 wkt2=-5.3368725e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.508574e-007 wpclm=-2.3611051e-008 wr=1 wtvoff=0 wu0=-5.9339327e-009 wua1=2.5344044e-017 wua=1.9445519e-017 wub1=-1.1253962e-024 wub=-3.1744322e-025 wuc1=-9.8477906e-018 wuc=-1.6185636e-017 wute=-2.7452583e-008 wvoffcv=8.2971572e-008 wvth0=-2.7658345e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.11 nmos a0=1.0800597 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29635114 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.100643 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79290591 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31356294 kt1l=0 kt2=-0.017501421 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1132954 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040683961 ua1=1.6559664e-009 ua=-7.8609378e-010 ub1=-2.3243083e-018 ub=3.2061309e-018 uc1=-5.6e-011 uc=1.1070566e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.0573125 voffl=0 vsat=75000 vth0=0.71889441 w0=5e-007 wa0=9.2126199e-008 wags=-7.6882295e-009 wbeta0=-3.1548252e-007 wint=1e-008 wk1=-2.6511136e-009 wkt1=-3.5962356e-008 wkt2=-4.9708381e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.3255568e-007 wr=1 wtvoff=0 wu0=-6.2009548e-009 wua1=2.2269354e-017 wua=1.7086427e-017 wub1=-8.9223229e-025 wub=-4.0509016e-025 wuc=-2.4981444e-017 wvoffcv=7.2905625e-008 wvth0=-3.2343586e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.12 nmos a0=0.13372839 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.46825513 alpha0=2.6346295e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=2.53e-010 cgidl=0.5 cgsl=1.1e-010 cgso=2.53e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0032954546 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.96194091 k2=0.019191068 k3=0 k3b=0 keta=-0.12409156 kt1=-0.29257841 kt1l=0 kt2=-0.024617727 ku0=0 kvsat=0 kvth0=0 la0=-1.6334972e-008 lags=-6.8085644e-008 lalpha0=-2.8223522e-013 ldelta=3.4528409e-009 level=54 lint=0 lk1=-1.0430342e-007 lk2=-3.339933e-008 lketa=3.0741152e-008 lkt1=-7.1335693e-009 lkt2=7.0437954e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.2430227e-006 lpclm=-1.7008694e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=6.4153784e-010 lua=2.9527314e-016 lub1=4.8961284e-025 lub=-3.5612601e-025 luc1=4.7587744e-017 luc=-7.0348871e-017 lvoffcv=-1.0703807e-007 lvth0=-5.8511842e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.41363636 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.5411576e-013 pags=9.6123512e-013 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23454659 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pketa=1.9486253e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.045205295 ua1=1.675e-009 ua=-6.8558591e-010 ub1=-5.2160045e-018 ub=3.6641068e-018 uc1=-2.1358339e-010 uc=2.8527975e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.21284091 voffl=0 vsat=75000 vth0=0.82418523 w0=5e-007 wa0=-2.9925391e-007 wags=-1.866476e-006 wint=1e-008 wketa=-3.7837384e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.13 nmos a0=0.63315593 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.62032529 alpha0=6.7617464e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0013214286 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.017320476 k3=0 k3b=0 keta=-0.043632179 kt1=-0.31240086 kt1l=0 kt2=-0.022382143 ku0=0 kvsat=0 kvth0=0 la0=-2.7354015e-007 lags=-1.4640177e-007 lalpha0=-2.4077004e-012 ldelta=4.4694643e-009 level=54 lint=0 lk2=-3.2435975e-008 lketa=-1.0695428e-008 lkt1=3.0749914e-009 lkt2=-4.4694643e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=7.0823131e-008 lpdiblc2=9.4484475e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.6062299e-009 lua=4.409931e-016 lub1=-6.5924598e-025 lub=-2.2579734e-025 luc1=9.2875468e-018 lvoff=-8.6260661e-009 lvth0=-1.168318e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.063999357 pdiblc1=0.39 pdiblc2=0.00133635 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.037506864 ua1=1.675e-009 ua=-9.6853729e-010 ub1=-2.9852107e-018 ub=3.4110414e-018 uc1=-1.3921407e-010 uc=1.4868e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10391036 voffcv=0.005 voffl=0 vsat=75000 vth0=0.73325579 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.14 nmos a0=1.1833631 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26737957 alpha0=9.1059211e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.481134 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=1.23e-010 cgidl=0.5 cgsl=1.1e-010 cgso=1.23e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027238636 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79722801 k2=-0.0074202574 k3=0 k3b=0 keta=-0.020978796 kt1=-0.3181779 kt1l=0 kt2=-0.017344176 ku0=0 kvsat=0 kvth0=0 la0=-9.4204186e-007 lags=2.8242727e-007 lalpha0=-1.0482912e-010 lbeta0=-4.1275172e-006 ldelta=2.7655057e-009 level=54 lint=0 lk1=-4.5948877e-008 lk2=-2.3759842e-009 lketa=-3.8219289e-008 lkt1=1.0094096e-008 lkt2=-6.568076e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.3827528e-007 lpclm=-1.3238476e-007 lpdiblc2=1.7934304e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.7090825e-009 lua1=2.3230248e-017 lua=2.4723621e-016 lub1=-1.5403867e-024 lub=8.2550345e-026 luc1=-1.0449463e-016 luc=5.5973835e-017 lvoff=1.3343565e-008 lvoffcv=7.6051406e-008 lvth0=7.0105569e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1138068 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23124865 pdiblc1=0.39 pdiblc2=0.00063792557 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.039891348 ua1=1.6558805e-009 ua=-8.0906659e-010 ub1=-2.2599921e-018 ub=3.1572573e-018 uc1=-4.5566188e-011 uc=1.02611e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12199236 voffcv=-0.05759375 voffl=0 vsat=75000 vth0=0.71786999 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.model nmos_3p3.15 nmos a0=1.0893 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29558 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.069 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.1e-010 cgdo=2.53e-010 cgidl=0.5 cgsl=1.1e-010 cgso=2.53e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79264 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31717 kt1l=0 kt2=-0.018 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.4e-009 toxm=8e-009 toxp=8.4e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040062 ua1=1.6582e-009 ua=-7.8438e-010 ub1=-2.4138e-018 ub=3.1655e-018 uc1=-5.6e-011 uc=1.082e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.05 voffl=0 vsat=75000 vth0=0.71857 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.5e-008 xpart=0 xtis=3 xw=-1e-008
.subckt nplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 r_rsh0='rsh_nplus_u_m' r_dw=-5e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.36e-3 r_tc2=6.5e-7 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model np_junction d cj=0.00096797 level=2
d1 3 1 np_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends nplus_u_m1
.endl nmos_3p3_s

.lib nmos_3p3_fs
.subckt nmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.007148
.param par_k=0.007008
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b nplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b nplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b nmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model nmos_3p3.0 nmos a0=0.11206719 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.32050776 alpha0=2.627733e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=19.907557 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0038636364 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95223909 k2=0.052721915 k3=0 k3b=0 keta=-0.14660298 kt1=-0.45797555 kt1l=0 kt2=-0.024695 ku0=0 kvsat=0 kvth0=0 la0=-3.0583422e-009 lags=-1.3683815e-008 lalpha0=-2.876129e-013 lbeta0=1.2151841e-007 ldelta=3.0068182e-009 level=54 lint=0 lk1=-9.4486255e-008 lk2=-3.9622207e-008 lketa=3.6813935e-008 lkt1=4.0235308e-008 lkt2=1.20015e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-4.5110649e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.4287103e-009 lua=6.7054848e-016 lub1=2.7447418e-025 lub=-7.5166395e-025 luc1=-3.6983864e-018 luc=-5.8253799e-017 lute=8.8056818e-008 lvoff=3.7921347e-009 lvsat=-0.0026417045 lvth0=-3.6607582e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.7078752e-015 pags=-1.1953845e-014 palpha0=-1.3367465e-020 paramchk=1 pbeta0=8.5415114e-016 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.36959505 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=5.2733156e-015 pketa=-2.3745402e-015 pkt1=-8.4689085e-015 pkt2=-2.9041139e-016 ppclm=8.3834934e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-6.3741029e-016 pua=-1.3848566e-022 pub1=-5.6267206e-032 pub=9.0672414e-032 puc1=1.7937174e-024 puc=5.3308427e-024 pute=-4.2707557e-014 pvag=0 pvoff=-1.4541923e-015 pvsat=1.2812267e-009 pvth0=4.2707557e-016 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.023766155 ua1=1.675e-009 ua=-1.1188622e-009 ub1=-4.191221e-018 ub=3.341622e-018 uc1=-4.2302273e-011 uc=2.2389524e-010 ute=-1.5663149 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12625494 voffcv=0.005 voffl=0 vsat=97266.234 vth0=0.64635471 w0=5e-007 wa0=-6.3254637e-009 wags=4.8736973e-008 walpha0=4.9509131e-014 wbeta0=1.4348835e-007 wint=1e-008 wk2=-1.9530798e-008 wketa=8.2761628e-009 wkt1=3.2591386e-008 wkt2=1.0755977e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.2412267e-008 wr=1 wtvoff=0 wu0=4.7228328e-009 wua=2.6992935e-016 wub1=3.4262081e-025 wub=-4.17125e-025 wuc1=-6.6433977e-018 wuc=-3.333668e-017 wute=1.0491274e-007 wvoff=5.3858974e-009 wvsat=-0.00012912338 wvth0=-1.4783981e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.1 nmos a0=1.0806312 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.47491359 alpha0=6.5351125e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=22.62283 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0015 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.746507 k2=0.023469038 k3=0 k3b=0 keta=-0.028392375 kt1=-0.33934486 kt1l=0 kt2=-0.020325321 ku0=0 kvsat=0 kvth0=0 la0=-4.7765472e-007 lags=-8.9342671e-008 lalpha0=-2.2022289e-012 lbeta0=-1.2089656e-006 ldelta=4.165e-009 level=54 lint=0 lk1=6.32247e-009 lk2=-2.5288297e-008 lketa=-2.1109261e-008 lkt1=-1.7893733e-008 lkt2=-9.409925e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=9.5689239e-008 lpdiblc2=8.80481e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.5419574e-009 lua=7.5232737e-016 lub1=-4.0025352e-025 lub=-6.207519e-025 luc1=5.12295e-018 luc=9.9674311e-018 lvoff=-2.7639238e-009 lvsat=0.001561875 lvth0=-2.274447e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.4787741e-014 pags=-9.965144e-015 palpha0=1.8516415e-020 paramchk=1 pbeta0=2.4698413e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.082248339 pdiblc1=0.39 pdiblc2=0.0013741 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=-2.7446888e-015 pketa=5.4040719e-015 pkt1=8.6784603e-015 pkt2=2.5437886e-016 ppclm=-2.8898622e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.2313712e-015 pua=-2.995459e-023 pub1=8.2051973e-032 pub=-9.9142683e-032 puc1=-2.4846307e-024 puc=-1.2039633e-023 pvag=0 pvoff=3.2241042e-016 pvsat=2.0705256e-009 pvth0=-5.679156e-016 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.029657487 ua1=1.675e-009 ua=-1.2857579e-009 ub1=-2.8142257e-018 ub=3.0744545e-018 uc1=-6.0305e-011 uc=8.466824e-011 ute=-1.3866071 vbm=-3 version=4.5 vfbcv=-1 voff=-0.11287523 voffcv=0.005 voffl=0 vsat=88687.5 vth0=0.61806264 w0=5e-007 wa0=-5.3427231e-008 wags=4.4678399e-008 walpha0=-1.5560013e-014 wbeta0=-3.5881772e-007 wint=1e-008 wk2=-3.1675243e-009 wketa=-7.5985556e-009 wkt1=-2.4032443e-009 wkt2=-3.6219107e-011 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=4.5419115e-008 wr=1 wtvoff=0 wu0=9.0899306e-010 wua=4.8437374e-017 wub1=6.0336771e-026 wub=-2.974725e-026 wuc1=2.087925e-018 wuc=2.1132713e-018 wute=1.7754464e-008 wvoff=1.7601776e-009 wvsat=-0.0017399375 wvth0=-1.2753387e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.2 nmos a0=1.2236495 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.25812408 alpha0=7.4780689e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.201637 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027295455 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79588952 k2=0.0060240997 k3=0 k3b=0 keta=-0.019643215 kt1=-0.32862431 kt1l=0 kt2=-0.021116071 ku0=0 kvsat=0 kvth0=0 la0=-6.4784645e-007 lags=1.6863685e-007 lalpha0=-8.3414465e-011 lbeta0=-3.0877458e-006 ldelta=2.7018409e-009 level=54 lint=0 lk1=-5.2442732e-008 lk2=-4.5288209e-009 lketa=-3.1520762e-008 lkt1=-3.0651179e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=-3.1400457e-008 lpdiblc2=1.7521438e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.7345577e-009 lua=1.9286754e-016 lub1=-7.5229142e-025 lub=-2.2684367e-025 luc=-6.999336e-018 lvoff=1.3342993e-008 lvth0=-3.0036269e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-4.4036219e-014 pags=4.6367549e-014 palpha0=-9.2783067e-018 paramchk=1 pbeta0=-3.1995815e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.1890464 pdiblc1=0.39 pdiblc2=0.00064161023 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=2.6769992e-015 pketa=-2.8220597e-015 pkt1=1.4865822e-014 ppclm=4.8454232e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.4846634e-015 pua=2.0214448e-023 pub1=1.2630432e-031 pub=-1.1464767e-031 puc=1.4395718e-024 pvag=0 pvoff=-1.4870619e-016 pvth0=-3.7848123e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032410861 ua1=1.675e-009 ua=-8.1562356e-010 ub1=-2.5183956e-018 ub=2.7434392e-018 uc1=-5.6e-011 uc=9.8926027e-011 ute=-1.3866071 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12641046 voffcv=0.005 voffl=0 vsat=90000 vth0=0.6014737 w0=5e-007 wa0=4.40803e-009 wags=-2.659998e-009 walpha0=7.7968964e-012 wbeta0=1.1760436e-007 wint=1e-008 wk2=-7.7235646e-009 wketa=-6.8584002e-010 wkt1=-7.6027077e-009 wkt2=1.7754464e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.2728176e-009 wr=1 wtvoff=0 wu0=6.9614246e-010 wua=6.2785193e-018 wub1=2.3149925e-026 wub=-1.6717846e-026 wuc=-9.2137918e-018 wute=1.7754464e-008 wvoff=2.1560739e-009 wvth0=-1.0050112e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.3 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.27500464 alpha0=6.6430893e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.892554 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=0.0055707643 k3=0 k3b=0 keta=-0.022798446 kt1=-0.3316925 kt1l=0 kt2=-0.021116071 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.18590321 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032237232 ua1=1.675e-009 ua=-7.963175e-010 ub1=-2.5937e-018 ub=2.7207321e-018 uc1=-5.6e-011 uc=9.8225393e-011 ute=-1.3866071 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12507482 voffcv=0.005 voffl=0 vsat=90000 vth0=0.60117304 w0=5e-007 wags=1.9813982e-009 walpha0=6.868137e-012 wbeta0=8.5576518e-008 wint=1e-008 wk2=-7.4555967e-009 wketa=-9.6832848e-010 wkt1=-6.1146375e-009 wkt2=1.7754464e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=7.1230911e-009 wr=1 wtvoff=0 wu0=8.4475741e-010 wua=8.3019875e-018 wub1=3.5793e-026 wub=-2.8194089e-026 wuc=-9.0696905e-018 wute=1.7754464e-008 wvoff=2.1411884e-009 wvth0=-1.0428972e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.4 nmos a0=0.10671673 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.35387843 alpha0=2.6294657e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=20.979738 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0038636364 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95223909 k2=0.038660657 k3=0 k3b=0 keta=-0.12272005 kt1=-0.37648295 kt1l=0 kt2=-0.014808861 ku0=0 kvsat=0 kvth0=0 la0=-1.6137164e-009 lags=-1.1017368e-008 lalpha0=-2.6600418e-013 lbeta0=-8.5415114e-008 ldelta=3.0068182e-009 level=54 lint=0 lk1=-9.4486255e-008 lk2=-3.5825667e-008 lketa=2.8576826e-008 lkt1=1.5769644e-008 lkt2=-3.1561582e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-7.5885948e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=3.8067177e-009 lua=3.7738605e-016 lub1=2.3542184e-025 lub=-8.3236674e-026 luc=-3.2397203e-017 lvoff=-8.7450729e-009 lvsat=0.0040720909 lvth0=-3.9687122e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.0072317e-015 pags=-1.3247072e-014 palpha0=-2.3847691e-020 paramchk=1 pbeta0=1.0121691e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.45365742 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=3.4319939e-015 pketa=1.620458e-015 pkt1=3.3969382e-015 pkt2=1.8223981e-015 ppclm=2.3309514e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.357439e-016 pua=3.6981203e-024 pub1=-3.7326821e-032 pub=-2.3351482e-031 puc=-7.2096064e-024 pvag=0 pvoff=4.6263534e-015 pvsat=-1.9749641e-009 pvth0=1.9206526e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.033298195 ua1=1.675e-009 ua=-6.0169576e-010 ub1=-3.6418527e-018 ub=2.2763308e-018 uc1=-5.6e-011 uc=1.5632343e-010 ute=-1.4346429 vbm=-3 version=4.5 vfbcv=-1 voff=-0.079820841 voffcv=0.005 voffl=0 vsat=76839.61 vth0=0.66075684 w0=5e-007 wa0=-3.7304877e-009 wags=3.25522e-008 walpha0=4.8668758e-014 wbeta0=-3.7651952e-007 wint=1e-008 wk2=-1.2711088e-008 wketa=-3.3070572e-009 wkt1=-6.932527e-009 wkt2=-3.7191798e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.8357985e-008 wr=1 wtvoff=0 wu0=9.9793159e-011 wua=1.9103635e-017 wub1=7.6177186e-026 wub=9.954125e-026 wuc=-5.6435009e-019 wute=4.1051786e-008 wvoff=-1.7134642e-008 wvsat=0.009777789 wvth0=-2.1769016e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.5 nmos a0=0.9680546 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.4396228 alpha0=6.7781531e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.030477 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0015 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.76834994 k2=0.0078158961 k3=0 k3b=0 keta=-0.0440595 kt1=-0.40772797 kt1l=0 kt2=-0.031191964 ku0=0 kvsat=0 kvth0=0 la0=-4.2366927e-007 lags=-5.3032112e-008 lalpha0=-2.298861e-012 lbeta0=-1.102773e-007 ldelta=4.165e-009 level=54 lint=0 lk1=-4.3805685e-009 lk2=-2.0711735e-008 lketa=-9.966845e-009 lkt1=3.1079706e-008 lkt2=4.8715625e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=3.9557623e-008 lpdiblc2=8.80481e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.804274e-009 lua=6.4479186e-016 lub1=-1.7057876e-025 lub=-3.4825707e-025 luc1=3.0687684e-017 luc=4.0042012e-018 lvoff=1.1113945e-008 lvsat=-0.00404005 lvth0=-1.7189014e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.3952024e-015 pags=-2.7575765e-014 palpha0=6.5383015e-020 paramchk=1 pbeta0=-2.8587971e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.2180583 pdiblc1=0.39 pdiblc2=0.0013741 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=5.1909737e-015 pk2=-4.9643217e-015 pkt1=-1.5073657e-014 pkt2=-2.5647103e-015 ppclm=2.4333971e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.5085237e-016 pua=2.2200133e-023 pub1=-2.9340286e-032 pub=-2.3130267e-031 puc1=-1.4883527e-023 puc=-9.1474668e-024 pvag=0 pvoff=-6.4083562e-015 pvsat=4.7874593e-009 pvth0=-3.2623115e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.031262366 ua1=1.675e-009 ua=-1.1474219e-009 ub1=-2.8132801e-018 ub=2.8171887e-018 uc1=-1.1862793e-010 uc=8.2034846e-011 ute=-1.4346429 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12034945 voffcv=0.005 voffl=0 vsat=93395 vth0=0.61484234 w0=5e-007 wa0=1.172439e-009 wags=6.1794432e-008 walpha0=-1.3343472e-013 wbeta0=4.1347359e-007 wint=1e-008 wk1=-1.0593824e-008 wk2=4.4242495e-009 wkt1=3.0762566e-008 wkt2=5.2341027e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-2.0448715e-008 wr=1 wtvoff=0 wu0=1.3062678e-010 wua=-1.8655574e-017 wub1=5.9878135e-026 wub=9.5026674e-026 wuc1=3.0374545e-017 wuc=3.390467e-018 wute=4.1051786e-008 wvoff=5.3851733e-009 wvsat=-0.004023075 wvth0=-1.1191538e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.6 nmos a0=1.2327382 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.28395177 alpha0=9.0834879e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.03504 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027295455 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79415202 k2=-0.0057098764 k3=0 k3b=0 keta=-0.021057318 kt1=-0.33925459 kt1l=0 kt2=-0.021813326 ku0=0 kvsat=0 kvth0=0 la0=-7.3864278e-007 lags=1.3221642e-007 lalpha0=-1.0232637e-010 lbeta0=-3.6857066e-006 ldelta=2.7018409e-009 level=54 lint=0 lk1=-3.5085045e-008 lk2=-4.6160653e-009 lketa=-3.7339441e-008 lkt1=-5.0403614e-008 lkt2=-6.2890172e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=2.8621373e-008 lpdiblc2=1.7521438e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.4291291e-009 lua=2.1691469e-016 lub1=7.0670219e-025 lub=-6.3772226e-025 luc1=-4.9767852e-017 luc=-1.4541809e-017 lute=3.430373e-007 lvoff=1.3036382e-008 lvth0=1.3228117e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=6.4031457e-014 palpha0=-1.0603512e-019 paramchk=1 pbeta0=-2.9947156e-014 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.22724843 pdiblc1=0.39 pdiblc2=0.00064161023 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-8.4184784e-015 pk2=2.7193127e-015 pkt1=2.4445753e-014 pkt2=3.0501733e-015 ppclm=1.9343645e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.3365305e-015 pua=8.5515769e-024 pub1=-5.8130758e-031 pub=8.4628446e-032 puc1=2.4137408e-023 puc=5.0976715e-024 pute=-1.6637309e-013 pvag=0 pvth0=-1.1657208e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.03650052 ua1=1.675e-009 ua=-7.8786125e-010 ub1=-3.550491e-018 ub=3.0604368e-018 uc1=-5.1018233e-011 uc=9.7619729e-011 ute=-1.7229095 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12196494 voffcv=0.005 voffl=0 vsat=90000 vth0=0.58928172 w0=5e-007 wags=-1.5186427e-008 walpha0=1.0614126e-014 wbeta0=1.9840421e-007 wint=1e-008 wk1=8.4269053e-010 wk2=-2.0325861e-009 wkt1=-2.4470223e-009 wkt2=5.1571306e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.6255164e-008 wr=1 wtvoff=0 wu0=-1.287342e-009 wua=-7.1861991e-018 wub1=5.237162e-025 wub=-1.7046166e-025 wuc1=-2.416157e-018 wuc=-8.5802375e-018 wute=1.8086111e-007 wvth0=-4.137003e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.7 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29718664 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.6661 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=-0.006171945 k3=0 k3b=0 keta=-0.024795 kt1=-0.3443 kt1l=0 kt2=-0.022442857 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23011343 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.036357464 ua1=1.675e-009 ua=-7.6614807e-010 ub1=-3.47975e-018 ub=2.9966007e-018 uc1=-5.6e-011 uc=9.6164093e-011 ute=-1.6885714 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.005 voffl=0 vsat=90000 vth0=0.59060586 w0=5e-007 wags=-8.7768718e-009 wbeta0=1.954065e-007 wint=1e-008 wk2=-1.7603827e-009 wkt2=8.2103571e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.4318863e-008 wr=1 wtvoff=0 wu0=-1.1535552e-009 wua=-6.3301854e-018 wub1=4.6552725e-025 wub=-1.6199035e-025 wuc=-8.06996e-018 wute=1.6420714e-007 wvth0=-5.3038907e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.8 nmos a0=0.10356864 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.27282829 alpha0=2.5770972e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.140826 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0038636364 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.94377247 k2=0.011777641 k3=0 k3b=0 keta=-0.12210189 kt1=-0.28182405 kt1l=0 kt2=-0.025384429 ku0=0 kvsat=0 kvth0=0 la0=-7.6373182e-010 lags=3.0978636e-008 lalpha0=-2.4034362e-013 ldelta=3.0068182e-009 level=54 lint=0 lk1=-9.0337611e-008 lk2=-2.8567253e-008 lketa=2.8273926e-008 lkt1=-9.558142e-009 lkt2=9.1390428e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.2282169e-006 lpclm=-9.2361767e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.5943995e-010 lua=2.405174e-016 lub1=4.5632098e-025 lub=-3.1413979e-025 luc1=4.7020919e-017 luc=-6.4329084e-017 lvoff=6.518816e-010 lvoffcv=-1.0576312e-007 lvsat=-0.00032391632 lvth0=-5.2688923e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.50656508 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=-6.3012337e-014 palpha0=-5.4255458e-020 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.2039517 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-4.9161428e-015 pk2=-5.1692271e-015 pketa=1.9793943e-015 pkt1=3.3410365e-014 pkt2=-3.000626e-015 pnoff=-1.455437e-012 ppclm=-5.5670466e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=3.9862803e-015 pua=1.6588748e-022 pub1=-2.9909231e-031 pub=4.0105376e-032 puc1=-5.5719789e-023 puc=3.0629672e-023 pvag=0 pvoff=-6.5090378e-015 pvoffcv=1.253293e-013 pvsat=3.2343045e-009 pvth0=1.7327786e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.046917138 ua1=1.675e-009 ua=-6.4392181e-010 ub1=-5.3452175e-018 ub=3.7731784e-018 uc1=-2.2591814e-010 uc=2.8957392e-010 ute=-1.5701989 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12421225 voffcv=0.2208431 voffl=0 vsat=90661.054 vth0=0.69023545 w0=5e-007 wags=1.2859661e-007 walpha0=1.1072542e-013 wbeta0=-5.6740897e-007 wint=1e-008 wk1=1.0032944e-008 wk2=1.9145286e-008 wketa=-4.0395803e-009 wkt1=-1.1910332e-007 wkt2=8.8128685e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=2.9702796e-006 wpclm=2.775433e-007 wr=1 wtvoff=0 wu0=-1.6038654e-008 wua=6.9141509e-017 wub1=2.0946644e-024 wub=-1.6742232e-024 wuc1=2.0135299e-016 wuc=-1.5846619e-016 wute=2.0168565e-007 wvoff=3.5469172e-008 wvoffcv=-2.5577408e-007 wvsat=-0.0066006214 wvth0=-5.6701171e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.9 nmos a0=0.57552494 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.63099948 alpha0=6.66555e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.044222 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0015 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.016627153 k3=0 k3b=0 keta=-0.0440595 kt1=-0.30292054 kt1l=0 kt2=-0.021810866 ku0=0 kvsat=0 kvth0=0 la0=-2.3202232e-007 lags=-1.4452524e-007 lalpha0=-2.2436855e-012 lbeta0=4.7336172e-008 ldelta=4.165e-009 level=54 lint=0 lk2=-3.0943514e-008 lketa=-9.966845e-009 lkt1=7.7913898e-010 lkt2=-8.3714133e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=6.6793883e-008 lpdiblc2=8.80481e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.2633967e-009 lua=3.7694084e-016 lub1=-6.7075952e-025 lub=-1.6556982e-025 luc1=7.3792611e-018 luc=5.0028276e-019 lvoff=-9.8892719e-009 lvth0=-9.668011e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.2849684e-013 pags=8.0843597e-014 paramchk=1 pbeta0=-4.7265167e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.048788318 pdiblc1=0.39 pdiblc2=0.0013741 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=7.1603368e-015 pkt1=2.0832514e-014 pkt2=4.2001037e-015 ppclm=-7.9409961e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=2.9008716e-016 pua=3.3960359e-022 pub1=5.6337391e-031 pub=-4.4778706e-031 puc1=1.2736955e-023 puc=-4.9953234e-024 pvag=0 pvoff=1.8480456e-014 pvth0=-1.2174701e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.038541716 ua1=1.675e-009 ua=-9.2233701e-010 ub1=-3.0450532e-018 ub=3.4699744e-018 uc1=-1.450168e-010 uc=1.572691e-010 ute=-1.5701989 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10269969 voffcv=0.005 voffl=0 vsat=90000 vth0=0.60243767 w0=5e-007 wa0=4.6632009e-007 wags=-1.6498693e-007 wbeta0=3.9718628e-007 wint=1e-008 wk2=-6.0170898e-009 wkt1=-9.343424e-008 wkt2=-5.8824982e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.8013621e-007 wr=1 wtvoff=0 wu0=-8.4954031e-009 wua=-2.8538117e-016 wub1=3.3452927e-025 wub=-6.7852432e-025 wuc1=6.1645354e-017 wuc=-8.5762118e-017 wute=2.0168565e-007 wvoff=-1.5529795e-008 wvth0=3.5079858e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.10 nmos a0=1.1745182 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.2675321 alpha0=9.0843837e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.509036 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027295455 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79743934 k2=-0.007425139 k3=0 k3b=0 keta=-0.021057318 kt1=-0.31503813 kt1l=0 kt2=-0.01681628 ku0=0 kvsat=0 kvth0=0 la0=-9.448243e-007 lags=2.8800094e-007 lalpha0=-1.0241585e-010 lbeta0=-4.075793e-006 ldelta=2.7018409e-009 level=54 lint=0 lk1=-4.5254914e-008 lk2=-2.3212866e-009 lketa=-3.7339441e-008 lkt1=1.5199068e-008 lkt2=-6.7806996e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.5328342e-007 lpclm=-1.5280581e-007 lpdiblc2=1.7521438e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.9351498e-009 lua1=2.5751614e-017 lua=2.4388945e-016 lub1=-1.7366835e-024 lub=1.6776843e-025 luc1=-1.1187747e-016 luc=6.3428033e-017 lute=-2.7287058e-008 lvoff=1.3036382e-008 lvoffcv=8.430588e-008 lvth0=7.3148658e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1288096 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.4432511e-013 pags=-1.205732e-013 paramchk=1 pbeta0=4.3230522e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23332588 pdiblc1=0.39 pdiblc2=0.00064161023 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=3.632817e-015 pkt1=-5.3293425e-014 pkt2=3.632817e-015 pnoff=1.8164085e-013 ppclm=2.3433486e-013 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-2.65014e-015 pua1=-3.0515663e-023 pua=-2.3413506e-023 pub1=2.3141044e-030 pub=-8.6987803e-031 puc1=9.7737308e-023 puc=-8.7296592e-023 pute=2.7246128e-013 pvag=0 pvoffcv=-9.9902467e-014 pvth0=-4.6500058e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040498226 ua1=1.65336e-009 ua=-8.1052911e-010 ub1=-2.1493188e-018 ub=3.1898582e-018 uc1=-4.4801054e-011 uc=1.0438863e-010 ute=-1.5472686 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12196494 voffcv=-0.065845277 voffl=0 vsat=90000 vth0=0.58816635 w0=5e-007 wa0=6.8990718e-008 wags=4.2708771e-009 wbeta0=-3.632817e-007 wint=1e-008 wk1=-3.0527874e-009 wkt1=-3.1143535e-008 wkt2=-5.4057867e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.5263937e-007 wpclm=-2.3456943e-008 wr=1 wtvoff=0 wu0=-6.024624e-009 wua1=2.5643414e-017 wua=1.9675215e-017 wub1=-1.1366728e-024 wub=-3.2382603e-025 wuc1=-9.7835144e-018 wuc=-1.6601388e-017 wute=-2.7273401e-008 wvoffcv=8.3951653e-008 wvth0=-2.8152872e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.11 nmos a0=1.0799412 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29636102 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.101049 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79290932 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.3135167 kt1l=0 kt2=-0.017495028 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1134659 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040691935 ua1=1.6559377e-009 ua=-7.8611576e-010 ub1=-2.323161e-018 ub=3.2066518e-018 uc1=-5.6e-011 uc=1.1073779e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.05740625 voffl=0 vsat=90000 vth0=0.58889857 w0=5e-007 wa0=9.3447686e-008 wags=-7.7985119e-009 wbeta0=-3.200079e-007 wint=1e-008 wk1=-2.689142e-009 wkt1=-3.6478212e-008 wkt2=-5.0421413e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.344571e-007 wr=1 wtvoff=0 wu0=-6.2899032e-009 wua1=2.2588793e-017 wua=1.733152e-017 wub1=-9.0503075e-025 wub=-4.109009e-025 wuc=-2.5339785e-017 wvoffcv=7.3951406e-008 wvth0=-3.2807533e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.12 nmos a0=0.13104451 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.45707702 alpha0=2.5881864e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=2.185e-010 cgidl=0.5 cgsl=9.5e-011 cgso=2.185e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0038636364 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.94477727 k2=0.013695045 k3=0 k3b=0 keta=-0.11903243 kt1=-0.29375227 kt1l=0 kt2=-0.024501818 ku0=0 kvsat=0 kvth0=0 la0=-1.4226912e-008 lags=-5.9303239e-008 lalpha0=-2.4577732e-013 ldelta=3.0068182e-009 level=54 lint=0 lk1=-9.0829964e-008 lk2=-2.9084952e-008 lketa=2.6769891e-008 lkt1=-6.2120864e-009 lkt2=6.1339091e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.0824545e-006 lpclm=-1.4811586e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=5.5866682e-010 lua=2.5713106e-016 lub1=4.2636682e-025 lub=-3.1012323e-025 luc1=4.144057e-017 luc=-6.1261515e-017 lvoffcv=-9.3211364e-008 lvth0=-5.0953541e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.20909091 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.3442985e-013 pags=8.3845218e-013 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23174773 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pketa=1.6997185e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.045310864 ua1=1.675e-009 ua=-6.3699727e-010 ub1=-5.1354364e-018 ub=3.6055045e-018 uc1=-2.0575259e-010 uc=2.737035e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.19522727 voffl=0 vsat=90000 vth0=0.68455682 w0=5e-007 wa0=-2.7434664e-007 wags=-1.7111269e-006 wint=1e-008 wketa=-3.4688132e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.13 nmos a0=0.622227 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.614476 alpha0=6.66555e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0015 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.01602454 k3=0 k3b=0 keta=-0.0440595 kt1=-0.312278 kt1l=0 kt2=-0.0224 ku0=0 kvsat=0 kvth0=0 la0=-2.5490633e-007 lags=-1.3642874e-007 lalpha0=-2.2436855e-012 ldelta=4.165e-009 level=54 lint=0 lk2=-3.0226405e-008 lketa=-9.966845e-009 lkt1=2.86552e-009 lkt2=-4.165e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=6.599859e-008 lpdiblc2=8.80481e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.292449e-009 lua=4.1095222e-016 lub1=-6.143375e-025 lub=-2.104158e-025 luc1=8.65487e-018 lvoff=-8.03845e-009 lvth0=-1.088731e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.066829 pdiblc1=0.39 pdiblc2=0.0013741 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.0376909 ua1=1.675e-009 ua=-9.50918e-010 ub1=-3.01155e-018 ub=3.40202e-018 uc1=-1.38843e-010 uc=1.4868e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.104255 voffcv=0.005 voffl=0 vsat=90000 vth0=0.602789 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.14 nmos a0=1.1814276 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26795983 alpha0=9.0843837e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.472653 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=8.85e-011 cgidl=0.5 cgsl=9.5e-011 cgso=8.85e-011 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027295455 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.7971336 k2=-0.007425139 k3=0 k3b=0 keta=-0.021057318 kt1=-0.31815716 kt1l=0 kt2=-0.017357671 ku0=0 kvsat=0 kvth0=0 la0=-9.2035509e-007 lags=2.759255e-007 lalpha0=-1.0241585e-010 lbeta0=-4.0324976e-006 ldelta=2.7018409e-009 level=54 lint=0 lk1=-4.4891087e-008 lk2=-2.3212866e-009 lketa=-3.7339441e-008 lkt1=9.8617193e-009 lkt2=-6.4168722e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.3509204e-007 lpclm=-1.2933712e-007 lpdiblc2=1.7521438e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.6697377e-009 lua1=2.2695464e-017 lua=2.4154458e-016 lub1=-1.5049254e-024 lub=8.0649951e-026 luc1=-1.0208906e-016 luc=5.468526e-017 lvoff=1.3036382e-008 lvoffcv=7.4300625e-008 lvth0=6.8491667e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1135227 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23097666 pdiblc1=0.39 pdiblc2=0.00064161023 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.039894859 ua1=1.6559282e-009 ua=-8.0855864e-010 ub1=-2.2631568e-018 ub=3.1574269e-018 uc1=-4.5780875e-011 uc=1.02726e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12196494 voffcv=-0.0574375 voffl=0 vsat=90000 vth0=0.5878844 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.model nmos_3p3.15 nmos a0=1.0893 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29558 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.069 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=9.5e-011 cgdo=2.185e-010 cgidl=0.5 cgsl=9.5e-011 cgso=2.185e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79264 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31717 kt1l=0 kt2=-0.018 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=7.8e-009 toxm=8e-009 toxp=7.8e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040062 ua1=1.6582e-009 ua=-7.8438e-010 ub1=-2.4138e-018 ub=3.1655e-018 uc1=-5.6e-011 uc=1.082e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.05 voffl=0 vsat=90000 vth0=0.58857 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1e-008 xpart=0 xtis=3 xw=5e-009
.subckt nplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 r_rsh0='rsh_nplus_u_m' r_dw=-5e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.36e-3 r_tc2=6.5e-7 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model np_junction d cj=0.00096797 level=2
d1 3 1 np_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends nplus_u_m1
.endl nmos_3p3_fs

.lib nmos_3p3_sf
.subckt nmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.007148
.param par_k=0.007008
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b nplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b nplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b nmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model nmos_3p3.0 nmos a0=0.11186736 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.32766 alpha0=2.6763946e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=19.903605 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0034090909 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.96652273 k2=0.056667113 k3=0 k3b=0 keta=-0.1512997 kt1=-0.46065123 kt1l=0 kt2=-0.024763831 ku0=0 kvsat=0 kvth0=0 la0=-3.2269331e-009 lags=-1.6641391e-008 lalpha0=-3.2302945e-013 lbeta0=1.3594315e-007 ldelta=3.3613636e-009 level=54 lint=0 lk1=-1.0562749e-007 lk2=-4.3701293e-008 lketa=4.0887819e-008 lkt1=4.4027381e-008 lkt2=1.309011e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-4.9487196e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.8792474e-009 lua=7.3404439e-016 lub1=3.0051191e-025 lub=-8.3010051e-025 luc1=-3.9327954e-018 luc=-6.4523339e-017 lute=9.3637987e-008 lvoff=4.0757735e-009 lvsat=-0.0028091396 lvth0=-4.0876103e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.778677e-015 pags=-1.2449405e-014 palpha0=-1.3921628e-020 paramchk=1 pbeta0=8.8956088e-016 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.37854122 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=5.4919265e-015 pketa=-2.4729792e-015 pkt1=-8.8199961e-015 pkt2=-3.024507e-016 ppclm=8.73104e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-6.638348e-016 pua=-1.4422673e-022 pub1=-5.8599823e-032 pub=9.4431335e-032 puc1=1.8680778e-024 puc=5.5518384e-024 pute=-4.4478044e-014 pvag=0 pvoff=-1.5144774e-015 pvsat=1.3343413e-009 pvth0=4.4478044e-016 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.023581366 ua1=1.675e-009 ua=-1.1909754e-009 ub1=-4.197398e-018 ub=3.4119198e-018 uc1=-4.2438636e-011 uc=2.2926756e-010 ute=-1.5684253 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12626439 voffcv=0.005 voffl=0 vsat=86133.117 vth0=0.77039529 w0=5e-007 wa0=-6.1333689e-009 wags=4.7087182e-008 walpha0=4.8005613e-014 wbeta0=1.3355442e-007 wint=1e-008 wk2=-1.8937677e-008 wketa=8.0445414e-009 wkt1=3.1555052e-008 wkt2=1.0429334e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=1.9698751e-008 wr=1 wtvoff=0 wu0=4.4895909e-009 wua=2.7097128e-016 wub1=3.271121e-025 wub=-4.0136608e-025 wuc1=-6.4416477e-018 wuc=-3.1807431e-017 wute=1.0375203e-007 wvoff=5.2223358e-009 wvsat=-0.00030073052 wvth0=-1.3833002e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.1 nmos a0=1.0915554 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.48250605 alpha0=6.6090188e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=22.627356 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0013571429 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.74629014 k2=0.024027296 k3=0 k3b=0 keta=-0.028451232 kt1=-0.33900277 kt1l=0 kt2=-0.020297566 ku0=0 kvsat=0 kvth0=0 la0=-5.0286783e-007 lags=-9.5612876e-008 lalpha0=-2.3286678e-012 lbeta0=-1.2531695e-006 ldelta=4.4078571e-009 level=54 lint=0 lk1=6.6911271e-009 lk2=-2.7054986e-008 lketa=-2.1764897e-008 lkt1=-1.8013338e-008 lkt2=-9.6878403e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=1.0096118e-007 lpdiblc2=9.31821e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.7629382e-009 lua=7.930064e-016 lub1=-4.1485807e-025 lub=-6.6750038e-025 luc1=5.1571929e-018 luc=9.2670883e-018 lvoff=-2.8907672e-009 lvsat=0.0018733393 lvth0=-2.4131129e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.4438924e-014 pags=-9.8249129e-015 palpha0=1.8255849e-020 paramchk=1 pbeta0=2.4350853e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.083544401 pdiblc1=0.39 pdiblc2=0.0013439 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=-2.7060651e-015 pketa=5.3280249e-015 pkt1=8.5563355e-015 pkt2=2.507992e-016 ppclm=-2.8491956e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.2140431e-015 pua=-2.9533064e-023 pub1=8.0897323e-032 pub=-9.774753e-032 puc1=-2.4496666e-024 puc=-1.187021e-023 pvag=0 pvoff=3.1787341e-016 pvsat=2.0413888e-009 pvth0=-5.599238e-016 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.029691776 ua1=1.675e-009 ua=-1.3065872e-009 ub1=-2.7947117e-018 ub=3.0930961e-018 uc1=-6.0262143e-011 uc=8.4580446e-011 ute=-1.3848214 vbm=-3 version=4.5 vfbcv=-1 voff=-0.11260451 voffcv=0.005 voffl=0 vsat=76951.786 vth0=0.73756201 w0=5e-007 wa0=-5.0565226e-008 wags=4.194112e-008 walpha0=-1.5087478e-014 wbeta0=-3.4216904e-007 wint=1e-008 wk2=-2.8631843e-009 wketa=-7.2515451e-009 wkt1=-2.5161865e-009 wkt2=-4.1870281e-011 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=4.2405096e-008 wr=1 wtvoff=0 wu0=8.0747734e-010 wua=4.6081741e-017 wub1=5.3588288e-026 wub=-2.4544774e-026 wuc1=2.0245179e-018 wuc=2.3534472e-018 wute=1.6540179e-008 wvoff=1.6294911e-009 wvsat=-0.0016870982 wvth0=-1.1862994e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.2 nmos a0=1.2251902 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.25756499 alpha0=7.5706791e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.218715 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.002725 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79597775 k2=0.0052544426 k3=0 k3b=0 keta=-0.019658689 kt1=-0.32933993 kt1l=0 kt2=-0.021098214 ku0=0 kvsat=0 kvth0=0 la0=-6.6456596e-007 lags=1.7656581e-007 lalpha0=-8.5936972e-011 lbeta0=-3.1787135e-006 ldelta=2.75275e-009 level=54 lint=0 lk1=-5.3430878e-008 lk2=-4.3398333e-009 lketa=-3.2403874e-008 lkt1=-2.9705368e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=-2.7026844e-008 lpdiblc2=1.7851584e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.6151023e-009 lua=1.9857306e-016 lub1=-7.5352353e-025 lub=-2.4286628e-025 luc=-6.9837022e-018 lvoff=1.3579168e-008 lvth0=-3.4480652e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-4.1797436e-014 pags=4.4010242e-014 palpha0=-8.8066015e-018 paramchk=1 pbeta0=-3.0369161e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.18931963 pdiblc1=0.39 pdiblc2=0.0006386625 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=2.5409017e-015 pketa=-2.6785874e-015 pkt1=1.411005e-014 ppclm=4.5990839e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.4091837e-015 pua=1.9186754e-023 pub1=1.1988306e-031 pub=-1.0881903e-031 puc=1.3663846e-024 pvag=0 pvoff=-1.4114603e-016 pvth0=-3.5923941e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032483545 ua1=1.675e-009 ua=-8.1531997e-010 ub1=-2.5148229e-018 ub=2.7421588e-018 uc1=-5.6e-011 uc=9.8010851e-011 ute=-1.3848214 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12621602 voffcv=0.005 voffl=0 vsat=78500 vth0=0.72046857 w0=5e-007 wa0=4.1755681e-009 wags=-2.5507436e-009 walpha0=7.2781831e-012 wbeta0=1.1006248e-007 wint=1e-008 wk2=-7.1995204e-009 wketa=-6.345102e-010 wkt1=-7.1060329e-009 wkt2=1.6540179e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.0414302e-009 wr=1 wtvoff=0 wu0=6.462041e-010 wua=5.8174289e-018 wub1=2.136867e-026 wub=-1.5394771e-026 wuc=-8.5858868e-018 wute=1.6540179e-008 wvoff=2.008846e-009 wvth0=-9.3568204e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.3 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.27520393 alpha0=6.7121679e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.901161 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=0.0048208929 k3=0 k3b=0 keta=-0.022895839 kt1=-0.3323075 kt1l=0 kt2=-0.021098214 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.18661964 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032322196 ua1=1.675e-009 ua=-7.954825e-010 ub1=-2.5901e-018 ub=2.7178964e-018 uc1=-5.6e-011 uc=9.7313179e-011 ute=-1.3848214 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12485946 voffcv=0.005 voffl=0 vsat=78500 vth0=0.72012411 w0=5e-007 wags=1.8458839e-009 walpha0=6.3984027e-012 wbeta0=7.9723661e-008 wint=1e-008 wk2=-6.9456841e-009 wketa=-9.0210134e-010 wkt1=-5.6964375e-009 wkt2=1.6540179e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=6.6359196e-009 wr=1 wtvoff=0 wu0=7.869817e-010 wua=7.7341875e-018 wub1=3.3345e-026 wub=-2.6265804e-026 wuc=-8.4493848e-018 wute=1.6540179e-008 wvoff=1.9947455e-009 wvth0=-9.7157009e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.4 nmos a0=0.10689312 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.35614518 alpha0=2.6705875e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=20.985833 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0034090909 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.96652273 k2=0.043846284 k3=0 k3b=0 keta=-0.12710186 kt1=-0.37899643 kt1l=0 kt2=-0.014401245 ku0=0 kvsat=0 kvth0=0 la0=-1.7844039e-009 lags=-1.2574141e-008 lalpha0=-2.9783362e-013 lbeta0=-9.3517938e-008 ldelta=3.3613636e-009 level=54 lint=0 lk1=-1.0562749e-007 lk2=-3.9983252e-008 lketa=3.1977949e-008 lkt1=1.7695179e-008 lkt2=-3.492865e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-8.4380551e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.2490518e-009 lua=4.2195702e-016 lub1=2.6245527e-025 lub=-9.7593592e-026 luc=-3.6357518e-017 lvoff=-9.6862495e-009 lvsat=0.0045138312 lvth0=-4.4329423e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.0934756e-015 pags=-1.4381348e-014 palpha0=-2.5889643e-020 paramchk=1 pbeta0=1.0988358e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.46474849 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=3.7258573e-015 pketa=1.7592093e-015 pkt1=3.6878001e-015 pkt2=1.9784404e-015 ppclm=2.5305384e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.6449187e-016 pua=4.0147707e-024 pub1=-4.0522919e-032 pub=-2.5350945e-031 puc=-7.8269268e-024 pvag=0 pvoff=5.0224835e-015 pvsat=-2.1440698e-009 pvth0=2.0851079e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032725347 ua1=1.675e-009 ua=-6.5842313e-010 ub1=-3.6760182e-018 ub=2.29126e-018 uc1=-5.6e-011 uc=1.6123011e-010 ute=-1.4339286 vbm=-3 version=4.5 vfbcv=-1 voff=-0.07880914 voffcv=0.005 voffl=0 vsat=64899.351 vth0=0.78637258 w0=5e-007 wa0=-3.7706055e-009 wags=3.3556722e-008 walpha0=5.0764006e-014 wbeta0=-3.8050353e-007 wint=1e-008 wk2=-1.2847784e-008 wketa=-3.4494299e-009 wkt1=-7.2309805e-009 wkt2=-3.8792949e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-2.1249703e-008 wr=1 wtvoff=0 wu0=1.4619976e-010 wua=1.8008954e-017 wub1=7.9456704e-026 wub=1.3094736e-025 wuc=5.103582e-019 wute=3.9866071e-008 wvoff=-1.7318909e-008 wvsat=0.0097853084 wvth0=-2.1422215e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.5 nmos a0=0.98260745 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.44253343 alpha0=6.854642e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.041625 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0013571429 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.76831276 k2=0.0086062399 k3=0 k3b=0 keta=-0.043717643 kt1=-0.40824973 kt1l=0 kt2=-0.031266454 ku0=0 kvsat=0 kvth0=0 la0=-4.4839871e-007 lags=-5.6632149e-008 lalpha0=-2.4317014e-012 lbeta0=-1.219717e-007 ldelta=4.4078571e-009 level=54 lint=0 lk1=-4.5404077e-009 lk2=-2.201083e-008 lketa=-1.0548002e-008 lkt1=3.2614365e-008 lkt2=5.1083916e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=4.231228e-008 lpdiblc2=9.31821e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=5.0779459e-009 lua=6.8279785e-016 lub1=-1.8106533e-025 lub=-3.7282285e-025 luc1=3.2202986e-017 luc=4.0692393e-018 lvoff=1.1643984e-008 lvsat=-0.0041874643 lvth0=-1.8251362e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.4339074e-015 pags=-2.8340758e-014 palpha0=6.7196838e-020 paramchk=1 pbeta0=-2.9381044e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21633117 pdiblc1=0.39 pdiblc2=0.0013439 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=5.334979e-015 pk2=-5.1020394e-015 pkt1=-1.5491823e-014 pkt2=-2.6358592e-015 ppclm=2.5009032e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.6058554e-016 pua=2.2815997e-023 pub1=-3.0154229e-032 pub=-2.3771936e-031 puc1=-1.5296418e-023 puc=-9.4012312e-024 pvag=0 pvoff=-6.5861336e-015 pvsat=4.9202705e-009 pvth0=-3.3528129e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.031100065 ua1=1.675e-009 ua=-1.1698757e-009 ub1=-2.8063699e-018 ub=2.8309252e-018 uc1=-1.1914311e-010 uc=8.1961957e-011 ute=-1.4339286 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12063313 voffcv=0.005 voffl=0 vsat=81960.714 vth0=0.73523913 w0=5e-007 wa0=1.1850475e-009 wags=6.0928114e-008 walpha0=-1.3175851e-013 wbeta0=4.1105337e-007 wint=1e-008 wk1=-1.0460743e-008 wk2=4.4618175e-009 wkt1=3.0376124e-008 wkt2=5.1683514e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-2.0668622e-008 wr=1 wtvoff=0 wu0=1.3854029e-010 wua=-1.8856196e-017 wub1=5.912594e-026 wub=9.9986385e-026 wuc1=2.9992977e-017 wuc=3.5972295e-018 wute=3.9866071e-008 wvoff=5.4430856e-009 wvsat=-0.0040663393 wvth0=-1.0759625e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.6 nmos a0=1.2339809 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.28346322 alpha0=9.1007216e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.044693 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.002725 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79422595 k2=-0.0057375564 k3=0 k3b=0 keta=-0.0209945 kt1=-0.33921309 kt1l=0 kt2=-0.021793862 ku0=0 kvsat=0 kvth0=0 la0=-7.5256056e-007 lags=1.3584281e-007 lalpha0=-1.0425632e-010 lbeta0=-3.755685e-006 ldelta=2.75275e-009 level=54 lint=0 lk1=-3.5895368e-008 lk2=-4.6548363e-009 lketa=-3.8043005e-008 lkt1=-5.0919976e-008 lkt2=-6.3534453e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=2.9503581e-008 lpdiblc2=1.7851584e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.432364e-009 lua=2.2115348e-016 lub1=7.0971302e-025 lub=-6.4823822e-025 luc1=-5.0277701e-017 luc=-1.4725443e-017 lute=3.4655156e-007 lvoff=1.3282019e-008 lvth0=1.3270713e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=6.3353669e-014 palpha0=-1.0491271e-019 paramchk=1 pbeta0=-2.9630159e-014 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.22691687 pdiblc1=0.39 pdiblc2=0.0006386625 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-8.3293668e-015 pk2=2.6905281e-015 pkt1=2.4186989e-014 pkt2=3.0178865e-015 ppclm=1.9138888e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.322383e-015 pua=8.4610564e-024 pub1=-5.751543e-031 pub=8.3732633e-032 puc1=2.3881908e-023 puc=5.0437114e-024 pute=-1.6461199e-013 pvag=0 pvth0=-1.1533814e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.036480486 ua1=1.675e-009 ua=-7.8835147e-010 ub1=-3.5425504e-018 ub=3.0585412e-018 uc1=-5.0977253e-011 uc=9.7494752e-011 ute=-1.7203348 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12198688 voffcv=0.005 voffl=0 vsat=78500 vth0=0.70918783 w0=5e-007 wags=-1.4852404e-008 walpha0=1.048079e-014 wbeta0=1.9272256e-007 wint=1e-008 wk1=8.3210458e-010 wk2=-1.9783209e-009 wkt1=-2.4162826e-009 wkt2=4.9583426e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.5817263e-008 wr=1 wtvoff=0 wu0=-1.2523428e-009 wua=-6.9926086e-018 wub1=5.0953922e-025 wub=-1.6567642e-025 wuc1=-2.385805e-018 wuc=-8.3407396e-018 wute=1.7590904e-007 wvth0=-3.9984673e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.7 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29703393 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.6695 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=-0.006202575 k3=0 k3b=0 keta=-0.024795 kt1=-0.3443 kt1l=0 kt2=-0.022428571 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.22986429 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.036337393 ua1=1.675e-009 ua=-7.6625821e-010 ub1=-3.47165e-018 ub=2.9937821e-018 uc1=-5.6e-011 uc=9.6023679e-011 ute=-1.6857143 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.005 voffl=0 vsat=78500 vth0=0.71051357 w0=5e-007 wags=-8.5233661e-009 wbeta0=1.897625e-007 wint=1e-008 wk2=-1.7095369e-009 wkt2=7.9732143e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.3905286e-008 wr=1 wtvoff=0 wu0=-1.1202366e-009 wua=-6.1473482e-018 wub1=4.5208125e-025 wub=-1.5731152e-025 wuc=-7.8368723e-018 wute=1.5946429e-007 wvth0=-5.1506964e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.8 nmos a0=0.10368409 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26826194 alpha0=2.6135308e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.140347 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0034090909 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95743806 k2=0.016113039 k3=0 k3b=0 keta=-0.12637977 kt1=-0.28048406 kt1l=0 kt2=-0.025514754 ku0=0 kvsat=0 kvth0=0 la0=-8.5378636e-010 lags=3.4571911e-008 lalpha0=-2.6873472e-013 ldelta=3.3613636e-009 level=54 lint=0 lk1=-1.0099431e-007 lk2=-3.1940611e-008 lketa=3.1609683e-008 lkt1=-1.0653613e-008 lkt2=1.0188312e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.3716655e-006 lpclm=-1.0377847e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.8200638e-010 lua=2.6903445e-016 lub1=5.0984495e-025 lub=-3.5114332e-025 luc1=5.2512691e-017 luc=-7.1885433e-017 lvoff=7.2259769e-010 lvoffcv=-1.1811564e-007 lvsat=-0.00035905475 lvth0=-5.8885304e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.68954029 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=-6.977796e-014 palpha0=-6.0080856e-020 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.20558963 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-5.4439881e-015 pk2=-5.7242461e-015 pketa=2.1919215e-015 pkt1=3.699763e-014 pkt2=-3.3228026e-015 pnoff=-1.611707e-012 ppclm=-6.1647793e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=4.4142864e-015 pua=1.8369878e-022 pub1=-3.3120579e-031 pub=4.4411482e-032 puc1=-6.1702412e-023 puc=3.3918374e-023 pvag=0 pvoff=-7.2079119e-015 pvoffcv=1.3878588e-013 pvsat=3.5815711e-009 pvth0=1.9188267e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.046878971 ua1=1.675e-009 ua=-6.8024396e-010 ub1=-5.4123917e-018 ub=3.8192473e-018 uc1=-2.3284907e-010 uc=2.9916081e-010 ute=-1.5700284 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12427998 voffcv=0.2365993 voffl=0 vsat=79204.029 vth0=0.81815039 w0=5e-007 wags=1.3681953e-007 walpha0=1.178056e-013 wbeta0=-5.6205724e-007 wint=1e-008 wk1=1.0674487e-008 wk2=1.973878e-008 wketa=-4.2978854e-009 wkt1=-1.2298302e-007 wkt2=9.1790777e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=3.1602098e-006 wpclm=2.8326196e-007 wr=1 wtvoff=0 wu0=-1.6484308e-008 wua=4.3648431e-017 wub1=2.1196956e-024 wub=-1.6644377e-024 wuc1=2.0779766e-016 wuc=-1.6155822e-016 wute=1.9978338e-007 wvoff=3.6109333e-008 wvoffcv=-2.7212918e-007 wvsat=-0.0070226885 wvth0=-5.8761136e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.9 nmos a0=0.58388391 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.63581483 alpha0=6.7425071e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.042948 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0013571429 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.017683205 k3=0 k3b=0 keta=-0.043717643 kt1=-0.30302683 kt1l=0 kt2=-0.021787246 ku0=0 kvsat=0 kvth0=0 la0=-2.4575569e-007 lags=-1.5288006e-007 lalpha0=-2.3745126e-012 lbeta0=4.9673545e-008 ldelta=4.4078571e-009 level=54 lint=0 lk2=-3.2741396e-008 lketa=-1.0548002e-008 lkt1=8.4320304e-010 lkt2=-8.8219755e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=7.0681467e-008 lpdiblc2=9.31821e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.5122507e-009 lua=3.9922365e-016 lub1=-7.0936697e-025 lub=-1.7562456e-025 luc1=7.820931e-018 luc=5.249858e-019 lvoff=-1.0449376e-008 lvth0=-1.0242633e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.3953946e-013 pags=8.4750542e-014 paramchk=1 pbeta0=-4.9549361e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.046649798 pdiblc1=0.39 pdiblc2=0.0013439 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=7.5063759e-015 pkt1=2.1839292e-014 pkt2=4.403083e-015 ppclm=-8.3247623e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=3.0410627e-016 pua=3.5601568e-022 pub1=5.906002e-031 pub=-4.6942736e-031 puc1=1.3352496e-023 puc=-5.2367334e-024 pvag=0 pvoff=1.9373565e-014 pvth0=-1.276307e-014 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.038388296 ua1=1.675e-009 ua=-9.355169e-010 ub1=-3.0217801e-018 ub=3.4750928e-018 uc1=-1.4521817e-010 uc=1.571796e-010 ute=-1.5700284 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10237415 voffcv=0.005 voffl=0 vsat=78500 vth0=0.7227726 w0=5e-007 wa0=4.6968521e-007 wags=-1.6617753e-007 wbeta0=4.0949885e-007 wint=1e-008 wk2=-6.2036165e-009 wkt1=-9.3260785e-008 wkt2=-5.9697177e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.7870699e-007 wr=1 wtvoff=0 wu0=-8.4251315e-009 wua=-2.9422783e-016 wub1=3.1223288e-025 wub=-6.5691059e-025 wuc1=6.0631174e-017 wuc=-8.47835e-017 wute=1.9978338e-007 wvoff=-1.6011211e-008 wvth0=3.8885457e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.10 nmos a0=1.1761657 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26705136 alpha0=9.1016136e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.515585 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.002725 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79751289 k2=-0.0074212337 k3=0 k3b=0 keta=-0.0209945 kt1=-0.31508994 kt1l=0 kt2=-0.016809446 ku0=0 kvsat=0 kvth0=0 la0=-9.6241665e-007 lags=2.9332373e-007 lalpha0=-1.043456e-010 lbeta0=-4.1522184e-006 ldelta=2.75275e-009 level=54 lint=0 lk1=-4.6104496e-008 lk2=-2.3650252e-009 lketa=-3.8043005e-008 lkt1=1.5439565e-008 lkt2=-6.9053359e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.5601523e-007 lpclm=-1.5548326e-007 lpdiblc2=1.7851584e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.9693306e-009 lua1=2.6210559e-017 lua=2.4846474e-016 lub1=-1.7674141e-024 lub=1.7018056e-025 luc1=-1.1390135e-016 luc=6.4547999e-017 lute=-2.7566602e-008 lvoff=1.3282019e-008 lvoffcv=8.5808379e-008 lvth0=7.4486913e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1289382 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.4658091e-013 pags=-1.2168642e-013 paramchk=1 pbeta0=4.362966e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23356279 pdiblc1=0.39 pdiblc2=0.0006386625 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=3.666358e-015 pkt1=-5.3785472e-014 pkt2=3.666358e-015 pnoff=1.833179e-013 ppclm=2.3649842e-013 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-2.6746082e-015 pua1=-3.0797407e-023 pua=-2.3629677e-023 pub1=2.3354701e-030 pub=-8.7790942e-031 puc1=9.8639696e-023 puc=-8.8102583e-023 pute=2.7497685e-013 pvag=0 pvoffcv=-1.0082485e-013 pvth0=-4.6929382e-015 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040489883 ua1=1.6533384e-009 ua=-8.1092276e-010 ub1=-2.147361e-018 ub=3.1893035e-018 uc1=-4.4621244e-011 uc=1.0426802e-010 ute=-1.5472461 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12198688 voffcv=-0.065916016 voffl=0 vsat=78500 vth0=0.70815167 w0=5e-007 wa0=6.7932842e-008 wags=4.4315284e-009 wbeta0=-3.605757e-007 wint=1e-008 wk1=-3.0300479e-009 wkt1=-3.076098e-008 wkt2=-5.3608541e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.515024e-007 wpclm=-2.3626216e-008 wr=1 wtvoff=0 wu0=-5.9633841e-009 wua1=2.5452403e-017 wua=1.9528659e-017 wub1=-1.1298083e-024 wub=-3.193221e-025 wuc1=-9.8541155e-018 wuc=-1.6299327e-017 wute=-2.7470215e-008 wvoffcv=8.3326318e-008 wvth0=-2.7809847e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.11 nmos a0=1.0800202 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29635443 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.100778 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79290705 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31354753 kt1l=0 kt2=-0.01749929 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1133523 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040686619 ua1=1.6559568e-009 ua=-7.8610111e-010 ub1=-2.3239259e-018 ub=3.2063045e-018 uc1=-5.6e-011 uc=1.1071637e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.05734375 voffl=0 vsat=78500 vth0=0.7088958 w0=5e-007 wa0=9.25663e-008 wags=-7.7249574e-009 wbeta0=-3.1698963e-007 wint=1e-008 wk1=-2.6637784e-009 wkt1=-3.6134154e-008 wkt2=-4.9945845e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.3318892e-007 wr=1 wtvoff=0 wu0=-6.2305777e-009 wua1=2.2375739e-017 wua=1.7168052e-017 wub1=-8.9649462e-025 wub=-4.0702534e-025 wuc=-2.5100784e-017 wvoffcv=7.3253906e-008 wvth0=-3.2498097e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.12 nmos a0=0.13319227 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.46602357 alpha0=2.6253409e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=2.415e-010 cgidl=0.5 cgsl=1.05e-010 cgso=2.415e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0034090909 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95850818 k2=0.018091864 k3=0 k3b=0 keta=-0.12307965 kt1=-0.29281318 kt1l=0 kt2=-0.024594545 ku0=0 kvsat=0 kvth0=0 la0=-1.5902956e-008 lags=-6.6286522e-008 lalpha0=-2.7475786e-013 ldelta=3.3613636e-009 level=54 lint=0 lk1=-1.0154007e-007 lk2=-3.2514471e-008 lketa=2.9926622e-008 lkt1=-6.9445773e-009 lkt2=6.8571818e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.2100909e-006 lpclm=-1.6558077e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=6.2454136e-010 lua=2.8745037e-016 lub1=4.7664136e-025 lub=-3.4669104e-025 luc1=4.6326986e-017 luc=-6.8485095e-017 lvoffcv=-1.0420227e-007 lvth0=-5.6961668e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.37272727 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.5011547e-013 pags=9.3628492e-013 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23398682 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pketa=1.898046e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.045226409 ua1=1.675e-009 ua=-6.7586818e-010 ub1=-5.1998909e-018 ub=3.6523864e-018 uc1=-2.1201723e-010 uc=2.829645e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.20931818 voffl=0 vsat=78500 vth0=0.81225955 w0=5e-007 wa0=-2.9434406e-007 wags=-1.8358528e-006 wint=1e-008 wketa=-3.7216588e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.13 nmos a0=0.63097014 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.61915543 alpha0=6.7425071e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0013571429 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.017061289 k3=0 k3b=0 keta=-0.043717643 kt1=-0.31237629 kt1l=0 kt2=-0.022385714 ku0=0 kvsat=0 kvth0=0 la0=-2.6976967e-007 lags=-1.4438377e-007 lalpha0=-2.3745126e-012 ldelta=4.4078571e-009 level=54 lint=0 lk2=-3.1988877e-008 lketa=-1.0548002e-008 lkt1=3.0326057e-009 lkt2=-4.4078571e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=6.9846904e-008 lpdiblc2=9.31821e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.5427376e-009 lua=4.3491445e-016 lub1=-6.5015893e-025 lub=-2.2268494e-025 luc1=9.1595271e-018 lvoff=-8.5071643e-009 lvth0=-1.1522139e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.064565286 pdiblc1=0.39 pdiblc2=0.0013439 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.037543671 ua1=1.675e-009 ua=-9.6501343e-010 ub1=-2.9904786e-018 ub=3.4092371e-018 uc1=-1.3913986e-010 uc=1.4868e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10397929 voffcv=0.005 voffl=0 vsat=78500 vth0=0.72316243 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.14 nmos a0=1.182976 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26749563 alpha0=9.1016136e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.479438 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=1.115e-010 cgidl=0.5 cgsl=1.05e-010 cgso=1.115e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.002725 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79720913 k2=-0.0074212337 k3=0 k3b=0 keta=-0.0209945 kt1=-0.31817375 kt1l=0 kt2=-0.017346875 ku0=0 kvsat=0 kvth0=0 la0=-9.3769676e-007 lags=2.8112459e-007 lalpha0=-1.043456e-010 lbeta0=-4.1084794e-006 ldelta=2.75275e-009 level=54 lint=0 lk1=-4.5736941e-008 lk2=-2.3650252e-009 lketa=-3.8043005e-008 lkt1=1.0047538e-008 lkt2=-6.5377812e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.376375e-007 lpclm=-1.3177414e-007 lpdiblc2=1.7851584e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.7011995e-009 lua1=2.31231e-017 lua=2.4609585e-016 lub1=-1.5332818e-024 lub=8.2169587e-026 luc1=-1.0401266e-016 luc=5.571566e-017 lvoff=1.3282019e-008 lvoffcv=7.5700625e-008 lvth0=6.9782212e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.11375 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23119425 pdiblc1=0.39 pdiblc2=0.0006386625 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.03989205 ua1=1.65589e-009 ua=-8.08965e-010 ub1=-2.260625e-018 ub=3.1572912e-018 uc1=-4.5609125e-011 uc=1.02634e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12198688 voffcv=-0.0575625 voffl=0 vsat=78500 vth0=0.70787288 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.model nmos_3p3.15 nmos a0=1.0893 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29558 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.069 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1.05e-010 cgdo=2.415e-010 cgidl=0.5 cgsl=1.05e-010 cgso=2.415e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79264 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31717 kt1l=0 kt2=-0.018 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=530 rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe=8.2e-009 toxm=8e-009 toxp=8.2e-009 toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040062 ua1=1.6582e-009 ua=-7.8438e-010 ub1=-2.4138e-018 ub=3.1655e-018 uc1=-5.6e-011 uc=1.082e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.05 voffl=0 vsat=78500 vth0=0.70857 w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1e-008 xpart=0 xtis=3 xw=-5e-009
.subckt nplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 r_rsh0='rsh_nplus_u_m' r_dw=-5e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.36e-3 r_tc2=6.5e-7 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model np_junction d cj=0.00096797 level=2
d1 3 1 np_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends nplus_u_m1
.endl nmos_3p3_sf

.lib pmos_3p3_t
.subckt pmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.00666
.param par_k=0.002833
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b pplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b pplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b pmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model pmos_3p3.0 pmos a0=1.0272635 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19081247 alpha0=1.1485698e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=39.773597 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.86959286 k2=0.029351195 k3=0 k3b=0 keta=-0.066404636 kt1=-0.28373805 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.0434818e-007 lags=1.0492091e-007 lalpha0=-3.0054064e-012 lbeta0=-3.6237273e-006 level=54 lint=0 lk1=4.91e-009 lk2=-2.4890454e-008 lketa=8.2658182e-009 lkt1=-1.5974545e-008 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=7.0823636e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.4492727e-009 lua1=1.7181818e-016 lua=1.0386891e-015 lub1=-6.7359091e-025 lub=-1.4361909e-025 luc1=5.8570909e-017 luc=8.4861818e-018 lvoff=-1.6014546e-009 lvth0=-7.6827273e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.7370909e-015 pags=-1.2080073e-014 palpha0=6.39288e-020 paramchk=1 pbeta0=1.1827636e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.35627558 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-2.0974909e-014 pk2=3.4158327e-015 pketa=3.6614618e-015 pkt1=1.9400727e-015 ppclm=6.5406545e-015 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-5.2642909e-016 pua1=-8.9345454e-023 pua=-1.9180342e-022 pub1=1.4950473e-031 pub=1.3557818e-033 puc1=-1.4057018e-023 puc=-4.4743636e-024 pvag=0 pvoff=8.3275636e-016 pvth0=2.3570182e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0077071688 ua1=1.1563636e-009 ua=-2.4381818e-012 ub1=-2.100161e-018 ub=6.7035533e-019 uc1=-2.5418182e-010 uc=8.6801065e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094658091 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.7506174 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.1112467e-008 wags=-2.3219283e-008 walpha0=-1.0325417e-013 wbeta0=2.1005299e-007 wint=-1e-008 wk1=6.7137132e-008 wk2=-2.1522854e-008 wketa=-7.3229236e-009 wkt1=-1.1172031e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.9266005e-008 wtvoff=0 wu0=6.0892675e-010 wua1=1.7869091e-016 wua=3.3100364e-018 wub1=-1.4002317e-025 wub=-4.8420779e-027 wuc1=4.0843636e-017 wuc=-1.3364176e-017 wvoff=-1.6655127e-009 wvth0=4.2938493e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.1 pmos a0=1.1510659 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19022326 alpha0=7.5504633e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=42.422959 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.011648 k2=-0.018784 k3=0 k3b=0 keta=-0.0050909592 kt1=-0.30703735 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.6624939e-007 lags=1.0521551e-007 lalpha0=-3.5014873e-011 lbeta0=-4.9484082e-006 level=54 lint=0 lk1=-6.6117551e-008 lk2=-8.2285714e-010 lketa=-2.239102e-008 lkt1=-4.324898e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=1.2067592e-007 lpdiblc2=2.4533143e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.1587837e-009 lua=8.5199265e-016 lub1=-6.0410204e-025 lub=-3.5234082e-025 luc1=-3.0738122e-017 luc=5.8519641e-017 lvoff=1.2890571e-008 lvth0=8.0902041e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.6645518e-014 pags=-3.0616751e-014 palpha0=-2.3899709e-018 paramchk=1 pbeta0=8.5195102e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.25657102 pdiblc1=0.1484 pdiblc2=0.00024628714 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=2.1589126e-014 pk2=-6.084e-015 pketa=1.1021878e-015 pkt1=-1.6167967e-014 ppclm=-2.1505078e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-9.8910367e-017 pua=-1.6858315e-022 pub1=9.6045061e-032 pub=9.5112882e-032 puc1=3.2542237e-024 puc=-7.4630909e-024 pvag=0 pvth0=1.5205225e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010288147 ua1=1.5e-009 ua=3.7095469e-010 ub1=-2.2391388e-018 ub=1.0877988e-018 uc1=-7.5563755e-011 uc=-1.3265853e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12364214 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.78216327 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=3.8929322e-008 wags=1.3854074e-008 walpha0=4.8045453e-012 wbeta0=2.7621551e-007 wint=-1e-008 wk1=-1.7990939e-008 wk2=-2.5231886e-009 wketa=-2.2043755e-009 wkt1=2.5044049e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=8.5357469e-008 wtvoff=0 wu0=-2.4611069e-010 wua=-4.3130498e-017 wub1=-3.3103837e-026 wub=-1.9235628e-025 wuc1=6.2211526e-018 wuc=-7.386721e-018 wvth0=5.9668408e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.2 pmos a0=1.2626103 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.15731682 alpha0=0.0020588939 alpha1=0 at=12000 b0=0 b1=0 beta0=44.45026 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95493474 k2=-0.010993416 k3=0 k3b=0 keta=-0.00016272403 kt1=-0.26850506 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-4.001026e-007 lags=1.4470325e-007 lalpha0=-2.415082e-009 lbeta0=-7.3811688e-006 level=54 lint=0 lk1=1.9383117e-009 lk2=-1.0171558e-008 lketa=-2.8304903e-008 lkt1=-5.0563636e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4545454e-007 lpclm=4.2841558e-008 lpdiblc2=4.4675455e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=3.0025909e-009 lua=8.1926494e-016 lub1=3.3323377e-025 lub=-6.9161688e-026 luc1=-7.8734805e-017 luc=9.5515247e-017 lvoff=-1.8220325e-008 lvoffcv=-2.1818182e-007 lvth0=-9.5551948e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9454546 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=3.4170078e-014 pags=-1.4866597e-014 palpha0=-2.3332535e-017 paramchk=1 pbeta0=-6.7464935e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32143299 pdiblc1=0.1484 pdiblc2=7.8434545e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-3.6710649e-014 pk2=8.9552104e-015 pketa=2.6125948e-015 pkt1=2.6293091e-014 ppclm=7.4952935e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-6.5690182e-016 pua=-1.5714468e-022 pub1=-1.7328156e-031 pub=-4.1208312e-033 puc1=2.5455553e-023 puc=-1.8553586e-023 pvag=0 pvoff=-1.1894494e-015 pvth0=4.2667013e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0087516409 ua1=1.5e-009 ua=3.9822779e-010 ub1=-3.0202519e-018 ub=8.5181617e-019 uc1=-3.5566519e-011 uc=-4.4095525e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097716396 voffcv=0.021818182 voffl=0 vsat=94000 vth0=-0.76745877 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-3.4170078e-009 wags=7.2894545e-010 walpha0=2.2256682e-011 wbeta0=4.0343221e-007 wint=-1e-008 wk1=3.0592208e-008 wk2=-1.5055864e-008 wketa=-3.463048e-009 wkt1=-1.0340166e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=4.9757922e-009 wtvoff=0 wu0=2.1888218e-010 wua=-5.2662561e-017 wub1=1.9133501e-025 wub=-1.0966152e-025 wuc1=-1.2279955e-017 wuc=1.8553586e-018 wvoff=9.9120779e-010 wvth0=3.6783584e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.3 pmos a0=1.2226 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17178714 alpha0=0.0018173857 alpha1=0 at=12000 b0=0 b1=0 beta0=43.712143 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95512857 k2=-0.012010571 k3=0 k3b=0 keta=-0.0029932143 kt1=-0.27356143 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32571714 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0090519 ua1=1.5e-009 ua=4.8015429e-010 ub1=-2.9869286e-018 ub=8.449e-019 uc1=-4.344e-011 uc=-3.4544e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.099538429 voffcv=0 voffl=0 vsat=94000 vth0=-0.76841429 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-7.5771429e-010 walpha0=1.9923429e-011 wbeta0=3.9668571e-007 wint=-1e-008 wk1=2.6921143e-008 wk2=-1.4160343e-008 wketa=-3.2017886e-009 wkt1=-7.7108571e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=1.2471086e-008 wtvoff=0 wu0=1.53192e-010 wua=-6.8377029e-017 wub1=1.7400686e-025 wub=-1.100736e-025 wuc1=-9.7344e-018 wvoff=8.7226286e-010 wvth0=4.1050286e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.4 pmos a0=0.66833429 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20459958 alpha0=1.2079775e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=38.238696 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99870273 k2=0.014249873 k3=0 k3b=0 keta=-0.10490303 kt1=-0.33225761 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-1.03128e-007 lags=6.9689636e-008 lalpha0=-3.0255502e-012 lbeta0=-2.7152909e-006 level=54 lint=0 lk1=-3.5426364e-008 lk2=-2.0467636e-008 lketa=2.2143527e-008 lkt1=5.3309091e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=2.7248545e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.8372909e-009 lua1=-2.562e-016 lua=7.4813818e-016 lub1=-2.9730909e-026 lub=-3.0903909e-025 luc1=-3.4608e-017 luc=1.2453182e-017 lvth0=-2.1407273e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-5.5371585e-014 pags=6.2401891e-015 palpha0=7.4403585e-020 paramchk=1 pbeta0=-3.5411055e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3781492 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=1.1159673e-015 pketa=-3.5549469e-015 pkt1=-6.6438982e-015 ppclm=2.9199702e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-2.0819854e-016 pua1=1.33224e-022 pua=-4.0716945e-023 pub1=-1.8530247e-031 pub=8.7374182e-032 puc1=3.4396015e-023 puc=-6.5372036e-024 pvag=0 pvth0=-5.2482182e-016 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0091928468 ua1=2.0124e-009 ua=-8.0522078e-011 ub1=-2.8876353e-018 ub=1.748897e-018 uc1=6.432e-012 uc=8.6704408e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.7710094 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.9775566e-007 wags=-3.0388584e-008 walpha0=-4.121738e-013 wbeta0=1.0082017e-006 wint=-1e-008 wk2=-1.3670166e-008 wketa=1.2696239e-008 wkt1=1.4058139e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.7891728e-008 wtvoff=0 wu0=-1.6362577e-010 wua1=-2.66448e-016 wua=4.3913662e-017 wub1=2.6946346e-025 wub=-5.6568377e-025 wuc1=-9.4675549e-017 wuc=-1.3313914e-017 wvth0=1.4897689e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.5 pmos a0=1.3454526 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19226653 alpha0=0.000123026 alpha1=0 at=12000 b0=0 b1=0 beta0=43.366204 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.97705 k2=-0.026847376 k3=0 k3b=0 keta=-0.0016565918 kt1=-0.28366163 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-4.4168718e-007 lags=7.5856163e-008 lalpha0=-5.8498663e-011 lbeta0=-5.2790449e-006 level=54 lint=0 lk1=-2.46e-008 lk2=8.0987755e-011 lketa=-2.947969e-008 lkt1=-2.3764898e-008 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=-5.9909388e-008 lpdiblc2=2.4533143e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.5601469e-009 lua=5.7398498e-016 lub1=9.5240816e-026 lub=-7.120898e-026 luc1=1.8185143e-017 luc=5.1804544e-017 lvoff=1.2890571e-008 lvth0=-3.242449e-010 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.4582136e-014 pags=-1.5349891e-014 palpha0=9.8215995e-018 paramchk=1 pbeta0=2.571262e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.55246506 pdiblc1=0.1484 pdiblc2=0.00024628714 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-6.5539994e-015 pketa=4.7882958e-015 pkt1=-6.0591673e-015 ppclm=7.2399282e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-3.0761926e-016 pua=-2.4019161e-023 pub1=-2.6761322e-031 pub=-5.1075673e-032 puc1=-2.2185874e-023 puc=-3.9712404e-024 pvag=0 pvth0=5.8960359e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097471347 ua1=1.5e-009 ua=2.6778433e-010 ub1=-3.1375788e-018 ub=1.2732368e-018 uc1=-9.9154286e-011 uc=8.0016841e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12364214 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.77464237 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-6.215178e-008 wags=1.2791576e-008 walpha0=-1.9906566e-011 wbeta0=-2.1427184e-007 wint=-1e-008 wk2=1.6697667e-009 wketa=-3.9902465e-009 wkt1=1.2888678e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-6.8507432e-008 wtvoff=0 wu0=3.5215673e-011 wua=1.0518093e-017 wub1=4.3408496e-025 wub=-2.8878406e-025 wuc1=1.8488229e-017 wuc=-1.844584e-017 wvth0=2.0559739e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.6 pmos a0=1.1189871 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16561084 alpha0=0.002173683 alpha1=0 at=12000 b0=0 b1=0 beta0=44.354662 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0137659 k2=-0.027452061 k3=0 k3b=0 keta=-0.0068224318 kt1=-0.33774851 kt1l=0 kt2=-0.016947818 ku0=0 kvsat=0 kvth0=0 la0=-1.6992857e-007 lags=1.0784299e-007 lalpha0=-2.519287e-009 lbeta0=-6.4651948e-006 level=54 lint=0 lk1=-6.8659091e-008 lk2=8.0661039e-010 lketa=-2.3280682e-008 lkt1=4.1139351e-008 lkt2=4.6581818e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4545454e-007 lpclm=2.0841896e-007 lpdiblc2=4.4675455e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.5779454e-009 lua=4.1154156e-016 lub1=-5.5351558e-025 lub=5.7264156e-026 luc1=-4.9745455e-017 luc=6.0010667e-017 lvoff=-2.0507727e-008 lvoffcv=-2.1818182e-007 lvth0=-1.3737662e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9454546 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-8.5520416e-014 pags=4.3007377e-015 palpha0=3.0854085e-017 paramchk=1 pbeta0=-5.4377143e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3288581 pdiblc1=0.1484 pdiblc2=7.8434545e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=3.2465626e-015 pkt1=-2.1392462e-014 pkt2=-2.4222546e-015 ppclm=-1.1147314e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=8.3913818e-017 pua=5.487148e-023 pub1=2.878281e-031 pub=-6.986227e-032 puc1=1.0381091e-023 puc=-9.1205299e-026 pvag=0 pvth0=1.2358442e-017 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097323026 ua1=1.5e-009 ua=4.0315384e-010 ub1=-2.5969484e-018 ub=1.1661759e-018 uc1=-4.2545455e-011 uc=1.1632475e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.095810227 voffcv=0.021818182 voffl=0 vsat=94000 vth0=-0.77376777 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=7.1267013e-008 wags=-3.583948e-009 walpha0=-3.7433637e-011 wbeta0=4.5314286e-007 wint=-1e-008 wk2=-6.4973683e-009 wkt1=2.5666423e-008 wkt2=2.0185455e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.1147314e-009 wtvoff=0 wu0=-2.910619e-010 wua=-5.5224108e-017 wub1=-2.878281e-026 wub=-2.7312856e-025 wuc1=-8.6509091e-018 wuc=-2.1679203e-017 wvth0=6.9590384e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.7 pmos a0=1.1019943 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17639514 alpha0=0.0019217543 alpha1=0 at=12000 b0=0 b1=0 beta0=43.708143 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.0273714 k3=0 k3b=0 keta=-0.0091505 kt1=-0.33363457 kt1l=0 kt2=-0.016482 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0098900971 ua1=1.5e-009 ua=4.44308e-010 ub1=-2.6523e-018 ub=1.1719023e-018 uc1=-4.752e-011 uc=7.1643143e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0=-0.77390514 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=6.2714971e-008 wags=-3.1538743e-009 walpha0=-3.4348229e-011 wbeta0=3.9876571e-007 wint=-1e-008 wk2=-6.172712e-009 wkt1=2.3527177e-008 wkt2=1.77632e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wtvoff=0 wu0=-2.8267051e-010 wua=-4.973696e-017 wub=-2.8011479e-025 wuc1=-7.6128e-018 wuc=-2.1688323e-017 wvth0=6.9602743e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.8 pmos a0=0.8879706 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.3341873 alpha0=9.723125e-006 alpha1=0 at=12000 b0=0 b1=0 beta0=37.805966 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99870273 k2=-0.00067810868 k3=0 k3b=0 keta=-0.088919542 kt1=-0.29596713 kt1l=0 kt2=-0.020842369 ku0=0 kvsat=0 kvth0=0 la0=-1.4725376e-007 lags=-2.4436508e-009 lalpha0=-2.2830898e-012 lbeta0=-2.3737058e-006 level=54 lint=0 lk1=-3.5426364e-008 lk2=-1.7691446e-008 lketa=1.7668152e-008 lkt1=-8.3979897e-009 lkt2=2.1773833e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=5.0559583e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.7890915e-009 lua1=-1.5583996e-016 lua=6.3071157e-016 lub1=-1.2857843e-025 lub=3.2915171e-026 luc1=8.8928926e-019 luc=-7.439668e-018 lvth0=-8.7733719e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.5381528e-015 pags=9.42428e-014 palpha0=-8.3139811e-019 paramchk=1 pbeta0=-7.708444e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32482036 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-2.2709854e-015 pketa=1.9050111e-015 pkt1=4.2520201e-015 pkt2=-2.6564076e-015 ppclm=7.6023645e-016 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.493953e-016 pua1=1.078475e-023 pua=1.0254352e-022 pub1=-6.4708497e-032 pub=-3.2981002e-031 puc1=-8.9106783e-024 puc=1.7732073e-023 pvag=0 pvth0=7.5670046e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011352976 ua1=1.8116799e-009 ua=3.4788822e-010 ub1=-2.5843988e-018 ub=9.2772209e-019 uc1=-8.5778578e-011 uc=1.3375779e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.76226585 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-7.0200638e-008 wags=-1.884856e-007 walpha0=2.4629388e-012 wbeta0=1.5361323e-006 wint=-1e-008 wk2=4.5419708e-009 wketa=-6.803611e-009 wkt1=-3.0216242e-008 wkt2=9.4871699e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=8.2952909e-008 wtvoff=0 wu0=-2.7989835e-009 wua1=-2.1569499e-017 wua=-4.7874691e-016 wub1=-1.0048507e-025 wub=4.3614967e-025 wuc1=1.7821357e-017 wuc=-7.0719038e-017 wvth0=4.2305517e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.9 pmos a0=1.1782327 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20788505 alpha0=0.00011108151 alpha1=0 at=12000 b0=0 b1=0 beta0=43.187318 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.97705 k2=-0.030551827 k3=0 k3b=0 keta=-0.0066799724 kt1=-0.30269355 kt1l=0 kt2=-0.010621998 ku0=0 kvsat=0 kvth0=0 la0=-2.9238479e-007 lags=6.0707474e-008 lalpha0=-5.296228e-011 lbeta0=-5.0643818e-006 level=54 lint=0 lk1=-2.46e-008 lk2=-2.7545864e-009 lketa=-2.3451633e-008 lkt1=-5.0347792e-009 lkt2=-2.9328019e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.407763e-008 lpdiblc2=2.4533143e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.4020669e-009 lua=6.4174442e-016 lub1=-1.8989494e-025 lub=1.5676208e-026 luc1=-2.4594545e-017 luc=7.3318673e-017 lvoff=-1.787102e-009 lvth0=-7.1445584e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.0756678e-013 pags=3.1315103e-015 palpha0=3.0672131e-018 paramchk=1 pbeta0=-4.7627532e-015 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.37778426 pdiblc1=0.1484 pdiblc2=0.00024628714 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-3.0945989e-015 pketa=-2.5659333e-015 pkt1=-2.8909912e-014 pkt2=3.5780184e-015 ppclm=-3.006488e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.3347616e-015 pua=-1.0668567e-022 pub1=8.0252392e-032 pub=-1.570756e-031 puc1=3.0005345e-023 puc=-3.0218479e-023 pvag=0 pvoff=1.7906761e-014 pvth0=1.4216818e-014 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010127025 ua1=1.5e-009 ua=3.2582253e-010 ub1=-2.4617658e-018 ub=9.6220002e-019 uc1=-3.4810909e-011 uc=-2.7758895e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094286796 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.76552347 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.4185662e-007 wags=-6.2630205e-009 walpha0=-5.3342836e-012 wbeta0=3.968961e-009 wint=-1e-008 wk2=6.1891978e-009 wketa=2.1382778e-009 wkt1=3.6107623e-008 wkt2=-2.981682e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.4460314e-007 wtvoff=0 wu0=-4.282509e-010 wua=-6.0288518e-017 wub1=-3.9040685e-025 wub=9.0680837e-026 wuc1=-6.0010691e-017 wuc=2.5182066e-017 wvoff=-3.5813523e-008 wvth0=-9.069076e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.10 pmos a0=1.1832393 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16685819 alpha0=0.0021426891 alpha1=0 at=12000 b0=0 b1=0 beta0=44.161948 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0137659 k2=-0.036023042 k3=0 k3b=0 keta=-0.0068224318 kt1=-0.29670927 kt1l=0 kt2=-0.012757219 ku0=0 kvsat=0 kvth0=0 la0=-2.9839274e-007 lags=1.0993971e-007 lalpha0=-2.4908914e-009 lbeta0=-6.233938e-006 level=54 lint=0 lk1=-6.8659091e-008 lk2=3.8108709e-009 lketa=-2.3280682e-008 lkt1=-1.2215919e-008 lkt2=-3.7053719e-010 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4545454e-007 lpclm=6.5657665e-008 lpdiblc2=4.4675455e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.3166262e-009 lua1=1.2483595e-016 lua=2.315961e-016 lub1=4.4029649e-026 luc1=1.3542397e-017 luc=5.9935909e-017 lvoff=2.8431167e-009 lvoffcv=-2.1818182e-007 lvth0=-4.4690083e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9454546 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.1205867e-014 pags=1.7427347e-015 palpha0=-3.7885537e-018 paramchk=1 pbeta0=-8.2590471e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34313423 pdiblc1=0.1484 pdiblc2=7.8434545e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-4.1863519e-016 pkt1=4.3700967e-014 pkt2=3.7127826e-015 ppclm=1.6302147e-013 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=4.0272326e-016 pua1=-1.5229986e-022 pua=2.7440495e-022 pub1=-4.4117708e-031 puc1=-6.6830088e-023 pvag=0 pvoff=-2.848803e-014 pvth0=3.7885537e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011031559 ua1=1.39597e-009 ua=6.676128e-010 ub1=-2.656703e-018 ub=9.7526352e-019 uc1=-6.6591694e-011 uc=-1.6606591e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.098145312 voffcv=0.021818182 voffl=0 vsat=94000 vth0=-0.7677531 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-7.1205867e-009 wags=-5.1057076e-009 walpha0=3.7885537e-013 wbeta0=6.8825393e-007 wint=-1e-008 wk2=3.9592281e-009 wkt1=-2.4401443e-008 wkt2=-3.0939855e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=-1.6302147e-008 wtvoff=0 wu0=-1.8761549e-009 wua1=1.2691655e-016 wua=-3.7786403e-016 wub1=4.4117708e-026 wub=-4.0215498e-026 wuc1=2.0685503e-017 wvoff=2.848803e-009 wvth0=-3.7885537e-010 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.11 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17785216 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.538555 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035641955 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29793086 kt1l=0 kt2=-0.012794273 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011163222 ua1=1.4084536e-009 ua=6.9077241e-010 ub1=-2.6523e-018 ub=9.7526352e-019 uc1=-6.5237455e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0=-0.7682 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-4.9314341e-009 wbeta0=6.0566345e-007 wint=-1e-008 wk2=3.9173646e-009 wkt1=-2.0031346e-008 wkt2=-2.7227073e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wtvoff=0 wu0=-1.8358826e-009 wua1=1.1168656e-016 wua=-3.5042354e-016 wub=-4.0215498e-026 wuc1=1.4002494e-017 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.12 pmos a0=0.88096455 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.31537636 alpha0=9.9689273e-006 alpha1=0 at=12000 b0=0 b1=0 beta0=37.959273 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99870273 k2=-0.00022481818 k3=0 k3b=0 keta=-0.089598545 kt1=-0.29898273 kt1l=0 kt2=-0.019895546 ku0=0 kvsat=0 kvth0=0 la0=-1.4740727e-007 lags=6.9618182e-009 lalpha0=-2.3660636e-012 lbeta0=-2.4506364e-006 level=54 lint=0 lk1=-3.5426364e-008 lk2=-1.7918091e-008 lketa=1.7858273e-008 lkt1=-7.9736364e-009 lkt2=1.9122727e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=5.0635454e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.7741818e-009 lua1=-1.5476364e-016 lua=6.4094546e-016 lub1=-1.3503636e-025 luc=-5.67e-018 lvth0=-8.0181818e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.33309909 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011073636 ua1=1.8095273e-009 ua=3.0010909e-010 ub1=-2.5944273e-018 ub=9.7125e-019 uc1=-8.4e-011 uc=1.267e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.76184364 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.13 pmos a0=1.19239 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20726 alpha0=0.00011054914 alpha1=0 at=12000 b0=0 b1=0 beta0=43.187714 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.97705 k2=-0.029934143 k3=0 k3b=0 keta=-0.0064665714 kt1=-0.29909 kt1l=0 kt2=-0.010919571 ku0=0 kvsat=0 kvth0=0 la0=-3.0312e-007 lags=6.102e-008 lalpha0=-5.2656171e-011 lbeta0=-5.0648571e-006 level=54 lint=0 lk1=-2.46e-008 lk2=-3.0634286e-009 lketa=-2.3707714e-008 lkt1=-7.92e-009 lkt2=-2.5757143e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.1077143e-008 lpdiblc2=2.4533143e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.2688571e-009 lua=6.3109714e-016 lub1=-1.8188571e-025 luc1=-2.16e-017 luc=7.0302857e-017 lvth0=-5.7257143e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.39221571 pdiblc1=0.1484 pdiblc2=0.00024628714 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010084286 ua1=1.5e-009 ua=3.1980571e-010 ub1=-2.5007286e-018 ub=9.7125e-019 uc1=-4.08e-011 uc=-2.5245714e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.76642857 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.14 pmos a0=1.1825286 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16634864 alpha0=0.002142727 alpha1=0 at=12000 b0=0 b1=0 beta0=44.230636 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0137659 k2=-0.035627909 k3=0 k3b=0 keta=-0.0068224318 kt1=-0.29914454 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.9128636e-007 lags=1.1011364e-007 lalpha0=-2.4912696e-009 lbeta0=-6.3163636e-006 level=54 lint=0 lk1=-6.8659091e-008 lk2=3.7690909e-009 lketa=-2.3280682e-008 lkt1=-7.8545455e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4545454e-007 lpclm=8.1927273e-008 lpdiblc2=4.4675455e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.3568182e-009 lua1=1.0963636e-016 lua=2.5898182e-016 luc1=6.8727273e-018 luc=5.9935909e-017 lvoffcv=-2.1818182e-007 lvth0=-4.0909091e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9454546 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34150727 pdiblc1=0.1484 pdiblc2=7.8434545e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010844318 ua1=1.4086364e-009 ua=6.2990182e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.4527273e-011 uc=-1.6606591e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0.021818182 voffl=0 vsat=94000 vth0=-0.76779091 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.model pmos_3p3.15 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17736 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.599 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035251 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29993 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.9e-009 toxm=7.9e-009 toxp=7.9e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.01098 ua1=1.4196e-009 ua=6.558e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.384e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0=-0.7682 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=0 xpart=0 xtis=3 xw=0
.subckt pplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 par=1 r_rsh0='rsh_pplus_u_m' r_dw=2.75e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.375e-3 r_tc2=1e-6 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model pn_junction d cj=0.00094344 level=2
d1 1 3 pn_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends pplus_u_m1
.endl pmos_3p3_t

.lib pmos_3p3_f
.subckt pmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.00666
.param par_k=0.002833
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b pplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b pplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b pmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model pmos_3p3.0 pmos a0=1.0088763 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20174918 alpha0=1.1235927e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=39.445349 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.8647782 k2=0.028918855 k3=0 k3b=0 keta=-0.065134512 kt1=-0.28422543 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-1.9069135e-007 lags=9.8918351e-008 lalpha0=-2.8123501e-012 lbeta0=-3.3940359e-006 level=54 lint=0 lk1=6.1568267e-009 lk2=-2.3507638e-008 lketa=7.447618e-009 lkt1=-1.5068185e-008 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=6.5671827e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.3274457e-009 lua1=1.6719545e-016 lua=9.8467082e-016 lub1=-6.4044033e-025 lub=-1.3426634e-025 luc1=5.5767486e-017 luc=8.2624703e-018 lvoff=-1.5583678e-009 lvth0=-7.3534153e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.7146703e-015 pags=-1.198112e-014 palpha0=6.3405134e-020 paramchk=1 pbeta0=1.1730752e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.35995623 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-2.0803095e-014 pk2=3.3878523e-015 pketa=3.6314694e-015 pkt1=1.9241808e-015 ppclm=6.4870775e-015 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-5.221169e-016 pua1=-8.8613591e-023 pua=-1.9023228e-022 pub1=1.4828008e-031 pub=1.3446761e-033 puc1=-1.3941872e-023 puc=-4.4377124e-024 pvag=0 pvoff=8.2593493e-016 pvth0=2.3377109e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0078719299 ua1=1.1573864e-009 ua=8.7644416e-011 ub1=-2.1477044e-018 ub=6.5842379e-019 uc1=-2.5233764e-010 uc=8.863003e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094667623 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.67663617 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.154901e-008 wags=-2.5751203e-008 walpha0=-1.0380713e-013 wbeta0=2.3377646e-007 wint=-1e-008 wk1=6.9370633e-008 wk2=-2.2539936e-008 wketa=-7.4415355e-009 wkt1=-1.1684779e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=3.1666898e-008 wtvoff=0 wu0=5.9859026e-010 wua1=1.8158523e-016 wua=-1.3940377e-017 wub1=-1.3505708e-025 wub=-5.017448e-027 wuc1=4.2084409e-017 wuc=-1.4595908e-017 wvoff=-1.6924896e-009 wvth0=4.7732695e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.1 pmos a0=1.1426483 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19126654 alpha0=7.4423186e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=42.301722 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0117326 k2=-0.018588529 k3=0 k3b=0 keta=-0.0053639133 kt1=-0.30910467 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.5597206e-007 lags=1.0403388e-007 lalpha0=-3.3647732e-011 lbeta0=-4.787946e-006 level=54 lint=0 lk1=-6.5556919e-008 lk2=-3.2403549e-010 lketa=-2.1720434e-008 lkt1=-2.9271156e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=1.1826689e-007 lpdiblc2=2.3704904e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.1273211e-009 lua=8.3628161e-016 lub1=-5.9114366e-025 lub=-3.4780972e-025 luc1=-2.9952355e-017 luc=5.7121833e-017 lvoff=1.2455386e-008 lvth0=7.6993553e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.7075901e-014 pags=-3.1408371e-014 palpha0=-2.4517655e-018 paramchk=1 pbeta0=8.7397887e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.25217946 pdiblc1=0.1484 pdiblc2=0.00025119377 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=2.214733e-014 pk2=-6.2413065e-015 pketa=1.1306857e-015 pkt1=-1.6586003e-014 ppclm=-2.2061108e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.0146777e-016 pua=-1.72942e-022 pub1=9.852838e-032 pub=9.7572098e-032 puc1=3.3383641e-024 puc=-7.6560549e-024 pvag=0 pvth0=1.5598367e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010331202 ua1=1.5e-009 ua=3.9172068e-010 ub1=-2.2487222e-018 ub=1.0960127e-018 uc1=-7.6682222e-011 uc=-1.1491615e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12338433 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.70748201 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=4.0977761e-008 wags=1.4058737e-008 walpha0=5.050231e-012 wbeta0=2.9506668e-007 wint=-1e-008 wk1=-1.8642534e-008 wk2=-2.8080536e-009 wketa=-2.3169788e-009 wkt1=2.6245925e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=9.0167278e-008 wtvoff=0 wu0=-2.6339567e-010 wua=-4.9371285e-017 wub1=-3.3106883e-026 wub=-2.0220479e-025 wuc1=6.6740899e-018 wuc=-8.0009433e-018 wvth0=6.367274e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.2 pmos a0=1.2624812 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.1574043 alpha0=0.0020546973 alpha1=0 at=12000 b0=0 b1=0 beta0=44.410558 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95248832 k2=-0.0097979054 k3=0 k3b=0 keta=8.6249554e-005 kt1=-0.2677292 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-3.983336e-007 lags=1.4426221e-007 lalpha0=-2.3862134e-009 lbeta0=-7.2932429e-006 level=54 lint=0 lk1=4.8252741e-009 lk2=-1.0767296e-008 lketa=-2.8195228e-008 lkt1=-5.2081178e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.39352e-007 lpclm=3.6423596e-008 lpdiblc2=4.4175626e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=3.0210454e-009 lua=8.2254984e-016 lub1=3.4323494e-025 lub=-6.8061407e-026 luc1=-7.9870808e-017 luc=9.5916655e-017 lvoff=-1.7922234e-008 lvoffcv=-2.157408e-007 lvth0=-9.7863494e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.946 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=3.5872446e-014 pags=-1.5607258e-014 palpha0=-2.4494972e-017 paramchk=1 pbeta0=-7.0826067e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32107112 pdiblc1=0.1484 pdiblc2=7.88813e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-3.853959e-014 pk2=9.4013629e-015 pketa=2.7427554e-015 pkt1=2.7603024e-014 ppclm=7.8687123e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-6.8962895e-016 pua=-1.6497369e-022 pub1=-1.8191452e-031 pub=-4.3261328e-033 puc1=2.672376e-023 puc=-1.9477934e-023 pvag=0 pvoff=-1.2487082e-015 pvth0=4.4792702e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0087371575 ua1=1.5e-009 ua=4.0327941e-010 ub1=-3.0352362e-018 ub=8.6053432e-019 uc1=-3.4663323e-011 uc=-4.4147189e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097813945 voffcv=0.0216 voffl=0 vsat=94000 vth0=-0.6927634 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-3.5915545e-009 wags=7.5813661e-010 walpha0=2.3605119e-011 wbeta0=4.2825183e-007 wint=-1e-008 wk1=3.2440732e-008 wk2=-1.5975284e-008 wketa=-3.6739399e-009 wkt1=-1.0950226e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=5.3623696e-009 wtvoff=0 wu0=2.316895e-010 wua=-5.6078614e-017 wub1=2.0295616e-025 wub=-1.1643187e-025 wuc1=-1.3010587e-017 wuc=1.9501336e-018 wvoff=1.0511012e-009 wvth0=3.9098384e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.3 pmos a0=1.2226 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17184786 alpha0=0.0018157893 alpha1=0 at=12000 b0=0 b1=0 beta0=43.680357 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95297143 k2=-0.010875929 k3=0 k3b=0 keta=-0.0027366607 kt1=-0.27294357 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32471786 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.009039625 ua1=1.5e-009 ua=4.8563321e-010 ub1=-3.0008714e-018 ub=8.5372e-019 uc1=-4.266e-011 uc=-3.4544e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.099608321 voffcv=0 voffl=0 vsat=94000 vth0=-0.69374321 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-8.0446429e-010 walpha0=2.1152679e-011 wbeta0=4.2116071e-007 wint=-1e-008 wk1=2.8582143e-008 wk2=-1.5034018e-008 wketa=-3.3993348e-009 wkt1=-8.1866071e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=1.3240536e-008 wtvoff=0 wu0=1.6264375e-010 wua=-7.2595804e-017 wub1=1.8474286e-025 wub=-1.16865e-025 wuc1=-1.0335e-017 wvoff=9.2608036e-010 wvth0=4.3583036e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.4 pmos a0=0.65645235 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.21104356 alpha0=1.1826838e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=37.990543 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99566618 k2=0.012709478 k3=0 k3b=0 keta=-0.10320034 kt1=-0.33242454 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-9.5523869e-008 lags=6.5010179e-008 lalpha0=-2.8274782e-012 lbeta0=-2.5313328e-006 level=54 lint=0 lk1=-3.3094297e-008 lk2=-1.9136714e-008 lketa=2.0738198e-008 lkt1=5.9583152e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=2.5024839e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.7194104e-009 lua1=-2.4129648e-016 lua=6.9948888e-016 lub1=-2.5045136e-026 lub=-2.899821e-025 luc1=-3.2836296e-017 luc=1.1729669e-017 lvth0=-1.9920781e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-5.3153436e-014 pags=5.9902112e-015 palpha0=7.1423027e-020 paramchk=1 pbeta0=-3.3992511e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.38016331 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=1.0712624e-015 pketa=-3.4125381e-015 pkt1=-6.377748e-015 ppclm=2.8029981e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.9985825e-016 pua1=1.2788713e-022 pua=-3.9085851e-023 pub1=-1.7787938e-031 pub=8.387403e-032 puc1=3.3018133e-023 puc=-6.2753276e-024 pvag=0 pvth0=-5.037978e-016 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0093531893 ua1=1.99446e-009 ua=-1.7033143e-011 ub1=-2.8941809e-018 ub=1.7312067e-018 uc1=4.9114909e-012 uc=8.7990522e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.69642702 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.9833372e-007 wags=-3.0677229e-008 walpha0=-4.1699029e-013 wbeta0=1.0048234e-006 wint=-1e-008 wk2=-1.3948967e-008 wketa=1.2733351e-008 wkt1=1.3860749e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=2.0957146e-008 wtvoff=0 wu0=-1.8647726e-010 wua1=-2.620638e-016 wua=4.1538729e-017 wub1=2.6057544e-025 wub=-5.7359242e-025 wuc1=-9.4257628e-017 wuc=-1.4256968e-017 wvth0=1.5262418e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.5 pmos a0=1.3375751 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19358686 alpha0=0.00012216672 alpha1=0 at=12000 b0=0 b1=0 beta0=43.26392 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.976558 k2=-0.02687001 k3=0 k3b=0 keta=-0.0021847972 kt1=-0.28433818 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-4.2791177e-007 lags=7.352905e-008 lalpha0=-5.6673338e-011 lbeta0=-5.1047406e-006 level=54 lint=0 lk1=-2.3769504e-008 lk2=1.7807606e-010 lketa=-2.8557385e-008 lkt1=-2.2870309e-008 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=-5.8989544e-008 lpdiblc2=2.3704904e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.5121617e-009 lua=5.5497308e-016 lub1=9.6101442e-026 lub=-6.8027043e-026 luc1=1.790912e-017 luc=5.0116107e-017 lvoff=1.2455386e-008 lvth0=-4.0309955e-010 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.4052143e-014 pags=-1.5240812e-014 palpha0=9.7518057e-018 paramchk=1 pbeta0=2.5529903e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.55232393 pdiblc1=0.1484 pdiblc2=0.00025119377 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-6.5074256e-015 pketa=4.7542695e-015 pkt1=-6.01611e-015 ppclm=7.1884801e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-3.0543328e-016 pua=-2.3848477e-023 pub1=-2.6571152e-031 pub=-5.0712722e-032 puc1=-2.2028218e-023 puc=-3.9430202e-024 pvag=0 pvth0=5.8541378e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097778795 ua1=1.5e-009 ua=2.791058e-010 ub1=-3.142432e-018 ub=1.2763808e-018 uc1=-9.9075017e-011 uc=9.3297873e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12338433 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.69968312 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-6.2333454e-008 wags=1.2828966e-008 walpha0=-2.025384e-011 wbeta0=-2.1489817e-007 wint=-1e-008 wk2=1.5811316e-009 wketa=-4.0019103e-009 wkt1=1.3119687e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-6.8909289e-008 wtvoff=0 wu0=2.9865002e-011 wua=1.0314601e-017 wub1=4.4055934e-025 wub=-2.9779989e-025 wuc1=1.8542271e-017 wuc=-1.9036287e-017 wvth0=2.2338617e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.6 pmos a0=1.1176952 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16577511 alpha0=0.0021717533 alpha1=0 at=12000 b0=0 b1=0 beta0=44.341063 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0136972 k2=-0.027348888 k3=0 k3b=0 keta=-0.0068457125 kt1=-0.33811161 kt1l=0 kt2=-0.01697494 ku0=0 kvsat=0 kvth0=0 la0=-1.6669444e-007 lags=1.0656941e-007 lalpha0=-2.4915822e-009 lbeta0=-6.3843867e-006 level=54 lint=0 lk1=-6.7890933e-008 lk2=7.4698326e-010 lketa=-2.3020218e-008 lkt1=4.1012519e-008 lkt2=4.6438207e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.39352e-007 lpclm=2.0626092e-007 lpdiblc2=4.4175626e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.5589835e-009 lua=4.0608197e-016 lub1=-5.5180911e-025 lub=5.7712398e-026 luc1=-4.9350708e-017 luc=5.934069e-017 lvoff=-2.0278287e-008 lvoffcv=-2.157408e-007 lvth0=-1.3585892e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.946 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-8.6896311e-014 pags=4.3699301e-015 palpha0=3.1350481e-017 paramchk=1 pbeta0=-5.5251989e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32904913 pdiblc1=0.1484 pdiblc2=7.88813e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=3.2987949e-015 pkt1=-2.1736635e-014 pkt2=-2.461225e-015 ppclm=-1.1326658e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=8.5263865e-017 pua=5.575428e-023 pub1=2.9245883e-031 pub=-7.0986249e-032 puc1=1.0548107e-023 puc=-9.2672655e-026 pvag=0 pvth0=1.255727e-017 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097384672 ua1=1.5e-009 ua=4.0443501e-010 ub1=-2.5970528e-018 ub=1.1705395e-018 uc1=-4.2459e-011 uc=1.5649873e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.095830735 voffcv=0.0216 voffl=0 vsat=94000 vth0=-0.69887884 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=7.3145043e-008 wags=-3.6783923e-009 walpha0=-3.8434543e-011 wbeta0=4.6508409e-007 wint=-1e-008 wk2=-6.6732628e-009 wkt1=2.6352452e-008 wkt2=2.0717382e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.1340266e-009 wtvoff=0 wu0=-2.9900464e-010 wua=-5.6691087e-017 wub1=-2.928102e-026 wub=-2.8073464e-025 wuc1=-8.878878e-018 wuc=-2.227732e-017 wvth0=7.151017e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.7 pmos a0=1.1010057 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17644486 alpha0=0.0019222957 alpha1=0 at=12000 b0=0 b1=0 beta0=43.701857 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.0272741 k3=0 k3b=0 keta=-0.0091505 kt1=-0.33400543 kt1l=0 kt2=-0.01651 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0098945529 ua1=1.5e-009 ua=4.45092e-010 ub1=-2.6523e-018 ub=1.1763177e-018 uc1=-4.74e-011 uc=7.5061857e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0=-0.69901486 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=6.4444971e-008 wags=-3.2408743e-009 walpha0=-3.5295729e-011 wbeta0=4.0976571e-007 wint=-1e-008 wk2=-6.342987e-009 wkt1=2.4176177e-008 wkt2=1.82532e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wtvoff=0 wu0=-2.9046801e-010 wua=-5.110896e-017 wub=-2.8784179e-025 wuc1=-7.8228e-018 wuc=-2.2286598e-017 wvth0=7.1522743e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.8 pmos a0=0.87540638 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.33412543 alpha0=9.5254751e-006 alpha1=0 at=12000 b0=0 b1=0 beta0=37.601303 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99566618 k2=-0.0021980746 k3=0 k3b=0 keta=-0.087399697 kt1=-0.29666254 kt1l=0 kt2=-0.02066331 ku0=0 kvsat=0 kvth0=0 la0=-1.3755908e-007 lags=-2.3548078e-009 lalpha0=-2.1321619e-012 lbeta0=-2.2168591e-006 level=54 lint=0 lk1=-3.3094297e-008 lk2=-1.6525108e-008 lketa=1.6503627e-008 lkt1=-7.8484113e-009 lkt2=2.0360792e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=4.7230737e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.6714324e-009 lua1=-1.4558948e-016 lua=5.8911437e-016 lub1=-1.2006485e-025 lub=3.1000449e-026 luc1=8.3755803e-019 luc=-6.9634759e-018 lvth0=-8.201616e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.4501221e-015 pags=8.8849145e-014 palpha0=-7.8381597e-019 paramchk=1 pbeta0=-7.2672783e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32908612 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-2.1410135e-015 pketa=1.7959845e-015 pkt1=4.0086707e-015 pkt2=-2.5043775e-015 ppclm=7.1672699e-016 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.4084519e-016 pua1=1.0167522e-023 pua=9.6674803e-023 pub1=-6.1005134e-032 pub=-3.109345e-031 puc1=-8.400707e-024 puc=1.671724e-023 pvag=0 pvth0=7.1339337e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011508627 ua1=1.7983391e-009 ua=4.0233366e-010 ub1=-2.5953331e-018 ub=9.3020973e-019 uc1=-8.5716307e-011 uc=1.3317671e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.68802184 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-7.0979742e-008 wags=-1.8206792e-007 walpha0=2.4136865e-012 wbeta0=1.4835887e-006 wint=-1e-008 wk2=4.3873228e-009 wketa=-6.7014347e-009 wkt1=-3.0126506e-008 wkt2=9.344692e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=8.378208e-008 wtvoff=0 wu0=-2.8376654e-009 wua1=-2.0835087e-017 wua=-4.7428243e-016 wub1=-1.0700731e-025 wub=4.1163392e-025 wuc1=1.7214564e-017 wuc=-6.9835979e-017 wvth0=4.9240544e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.9 pmos a0=1.1722707 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20910427 alpha0=0.00011002657 alpha1=0 at=12000 b0=0 b1=0 beta0=43.086027 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.976558 k2=-0.030611931 k3=0 k3b=0 keta=-0.0071507123 kt1=-0.30282331 kt1l=0 kt2=-0.010678274 ku0=0 kvsat=0 kvth0=0 la0=-2.8242886e-007 lags=5.8655514e-008 lalpha0=-5.1176698e-011 lbeta0=-4.8934045e-006 level=54 lint=0 lk1=-2.3769504e-008 lk2=-2.6591455e-009 lketa=-2.2657878e-008 lkt1=-4.8419541e-009 lkt2=-2.8366187e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.3288533e-008 lpdiblc2=2.3704904e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.3220281e-009 lua=6.2016345e-016 lub1=-1.8354751e-025 lub=1.5271135e-026 luc1=-2.378795e-017 luc=7.086732e-017 lvoff=-1.7409232e-009 lvth0=-6.9145954e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.0489184e-013 pags=3.0536365e-015 palpha0=2.9909383e-018 paramchk=1 pbeta0=-4.6443141e-015 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.37814802 pdiblc1=0.1484 pdiblc2=0.00025119377 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-3.0176431e-015 pketa=-2.5021242e-015 pkt1=-2.8190987e-014 pkt2=3.489041e-015 ppclm=-2.9317233e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.301569e-015 pua=-1.0403264e-022 pub1=7.8256693e-032 pub=-1.5316948e-031 puc1=2.9259179e-023 puc=-2.9467012e-023 pvag=0 pvoff=1.746146e-014 pvth0=1.3863278e-014 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010175439 ua1=1.5e-009 ua=3.3870848e-010 ub1=-2.4652457e-018 ub=9.6244193e-019 uc1=-3.52542e-011 uc=-2.6312627e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094293534 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.69065918 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.4099098e-007 wags=-6.2574519e-009 walpha0=-5.3214657e-012 wbeta0=3.9093553e-009 wint=-1e-008 wk2=6.1836949e-009 wketa=2.1061652e-009 wkt1=3.5856399e-008 wkt2=-2.9369032e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.4532708e-007 wtvoff=0 wu0=-4.5913295e-010 wua=-6.2996698e-017 wub1=-3.9237991e-025 wub=8.8344941e-026 wuc1=-5.9957334e-017 wuc=2.4803882e-017 wvoff=-3.578168e-008 wvth0=-8.8655847e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.10 pmos a0=1.1829466 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.1669723 alpha0=0.002140198 alpha1=0 at=12000 b0=0 b1=0 beta0=44.155152 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0136972 k2=-0.036022469 k3=0 k3b=0 keta=-0.0068457125 kt1=-0.29670156 kt1l=0 kt2=-0.012755062 ku0=0 kvsat=0 kvth0=0 la0=-2.9511192e-007 lags=1.087083e-007 lalpha0=-2.4630203e-009 lbeta0=-6.1635247e-006 level=54 lint=0 lk1=-6.7890933e-008 lk2=3.7685735e-009 lketa=-2.3020218e-008 lkt1=-1.2114597e-008 lkt2=-3.6939483e-010 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.39352e-007 lpclm=6.4791222e-008 lpdiblc2=4.4175626e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.3015701e-009 lua1=1.2356248e-016 lua=2.2878304e-016 lub1=4.3893906e-026 luc1=1.3444942e-017 luc=5.9265346e-017 lvoff=2.8343515e-009 lvoffcv=-2.157408e-007 lvth0=-4.4220735e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.946 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.1057185e-014 pags=1.7390958e-015 palpha0=-3.780643e-018 paramchk=1 pbeta0=-8.2418018e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34321309 pdiblc1=0.1484 pdiblc2=7.88813e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-4.1776105e-016 pkt1=4.3609717e-014 pkt2=3.7050301e-015 ppclm=1.6268107e-013 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=4.0188235e-016 pua1=-1.5198185e-022 pua=2.7383197e-022 pub1=-4.4025588e-031 puc1=-6.6690543e-023 pvag=0 pvoff=-2.8428545e-014 pvth0=3.780643e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.01103441 ua1=1.3959912e-009 ua=6.6815328e-010 ub1=-2.6566947e-018 ub=9.7529642e-019 uc1=-6.6595019e-011 uc=-1.6546655e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.098144776 voffcv=0.0216 voffl=0 vsat=94000 vth0=-0.69275726 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-7.1142556e-009 wags=-5.1509361e-009 walpha0=3.7851852e-013 wbeta0=6.9375436e-007 wint=-1e-008 wk2=3.995242e-009 wkt1=-2.4581904e-008 wkt2=-3.1187122e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=-1.6287652e-008 wtvoff=0 wu0=-1.8930146e-009 wua1=1.2793085e-016 wua=-3.8106455e-016 wub1=4.4078482e-026 wub=-4.0585597e-026 wuc1=2.0808425e-017 wvoff=2.84627e-009 wvth0=-3.7851852e-010 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.11 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17785619 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.538059 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035645159 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29791448 kt1l=0 kt2=-0.012792045 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011164724 ua1=1.4083623e-009 ua=6.9105907e-010 ub1=-2.6523e-018 ub=9.7529642e-019 uc1=-6.5248909e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0=-0.6932 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-4.9768176e-009 wbeta0=6.1123732e-007 wint=-1e-008 wk2=3.9534157e-009 wkt1=-2.0215693e-008 wkt2=-2.7477641e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wtvoff=0 wu0=-1.8527781e-009 wua1=1.1271441e-016 wua=-3.5364845e-016 wub=-4.0585597e-026 wuc1=1.4131358e-017 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.12 pmos a0=0.86832964 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.31597309 alpha0=9.7661218e-006 alpha1=0 at=12000 b0=0 b1=0 beta0=37.749218 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99566618 k2=-0.0017606545 k3=0 k3b=0 keta=-0.088067836 kt1=-0.29966618 kt1l=0 kt2=-0.019731636 ku0=0 kvsat=0 kvth0=0 la0=-1.3770366e-007 lags=6.5035316e-009 lalpha0=-2.2103091e-012 lbeta0=-2.2893145e-006 level=54 lint=0 lk1=-3.3094297e-008 lk2=-1.6738569e-008 lketa=1.6682688e-008 lkt1=-7.4487433e-009 lkt2=1.7863906e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=4.7302195e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.65739e-009 lua1=-1.4457577e-016 lua=5.9875293e-016 lub1=-1.2614711e-025 luc=-5.296752e-018 lvth0=-7.4903564e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.33743927 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011225709 ua1=1.7962618e-009 ua=3.5504727e-010 ub1=-2.6060018e-018 ub=9.7125e-019 uc1=-8.4e-011 uc=1.26214e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.68753091 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.13 pmos a0=1.1863276 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.2084804 alpha0=0.00010949602 alpha1=0 at=12000 b0=0 b1=0 beta0=43.086417 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.976558 k2=-0.029995411 k3=0 k3b=0 keta=-0.0069407257 kt1=-0.2992484 kt1l=0 kt2=-0.010971086 ku0=0 kvsat=0 kvth0=0 la0=-2.9288667e-007 lags=5.8959965e-008 lalpha0=-5.0878499e-011 lbeta0=-4.8938676e-006 level=54 lint=0 lk1=-2.3769504e-008 lk2=-2.9600072e-009 lketa=-2.2907342e-008 lkt1=-7.6526208e-009 lkt2=-2.4887582e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.0365578e-008 lpdiblc2=2.3704904e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.1922605e-009 lua=6.097913e-016 lub1=-1.7574525e-025 luc1=-2.0870784e-017 luc=6.7929433e-017 lvth0=-5.5324142e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.39263726 pdiblc1=0.1484 pdiblc2=0.00025119377 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010129663 ua1=1.5e-009 ua=3.3242766e-010 ub1=-2.5043663e-018 ub=9.7125e-019 uc1=-4.1232e-011 uc=-2.3839657e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.69154309 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.14 pmos a0=1.1822374 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16645875 alpha0=0.0021402357 alpha1=0 at=12000 b0=0 b1=0 beta0=44.22432 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0136972 k2=-0.03562414 k3=0 k3b=0 keta=-0.0068457125 kt1=-0.2991524 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.8802745e-007 lags=1.0888169e-007 lalpha0=-2.4633972e-009 lbeta0=-6.2456962e-006 level=54 lint=0 lk1=-6.7890933e-008 lk2=3.7269223e-009 lketa=-2.3020217e-008 lkt1=-7.7666688e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.39352e-007 lpclm=8.101067e-008 lpdiblc2=4.4175626e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.3416381e-009 lua1=1.0840975e-016 lua=2.5608433e-016 luc1=6.7958352e-018 luc=5.9265346e-017 lvoffcv=-2.157408e-007 lvth0=-4.04514e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.946 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3415892 pdiblc1=0.1484 pdiblc2=7.88813e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010845675 ua1=1.408746e-009 ua=6.301608e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.45204e-011 uc=-1.6546655e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0.0216 voffl=0 vsat=94000 vth0=-0.692795 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.model pmos_3p3.15 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17736 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.599 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.6e-011 cgdo=1.116e-010 cgidl=7.5 cgsl=3.6e-011 cgso=1.116e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035251 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29993 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.5e-009 toxm=7.9e-009 toxp=7.5e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.01098 ua1=1.4196e-009 ua=6.558e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.384e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0=-0.6932 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-1.2e-008 xpart=0 xtis=3 xw=1e-008
.subckt pplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 par=1 r_rsh0='rsh_pplus_u_m' r_dw=2.75e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.375e-3 r_tc2=1e-6 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model pn_junction d cj=0.00094344 level=2
d1 1 3 pn_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends pplus_u_m1
.endl pmos_3p3_f

.lib pmos_3p3_s
.subckt pmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.00666
.param par_k=0.002833
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b pplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b pplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b pmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model pmos_3p3.0 pmos a0=1.0456883 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.1800417 alpha0=1.1734592e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=40.100221 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.87469564 k2=0.029736614 k3=0 k3b=0 keta=-0.067725055 kt1=-0.28327733 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.1845471e-007 lags=1.1100987e-007 lalpha0=-3.2039603e-012 lbeta0=-3.8596059e-006 level=54 lint=0 lk1=3.4485427e-009 lk2=-2.6287876e-008 lketa=9.1402523e-009 lkt1=-1.6892981e-008 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=7.6191219e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.570498e-009 lua1=1.7583709e-016 lua=1.092789e-015 lub1=-7.0652532e-025 lub=-1.5325276e-025 luc1=6.134421e-017 luc=8.679411e-018 lvoff=-1.6389133e-009 lvth0=-8.0025899e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.7472452e-015 pags=-1.2124889e-014 palpha0=6.4165969e-020 paramchk=1 pbeta0=1.1871516e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3525051 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-2.1052724e-014 pk2=3.4285051e-015 pketa=3.6750454e-015 pkt1=1.9472702e-015 ppclm=6.5649197e-015 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-5.2838208e-016 pua1=-8.9676916e-023 pua=-1.9251499e-022 pub1=1.5005937e-031 pub=1.3608116e-033 puc1=-1.4109168e-023 puc=-4.490963e-024 pvag=0 pvoff=8.358458e-016 pvth0=2.3657625e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.007549639 ua1=1.1565682e-009 ua=-8.9886117e-011 ub1=-2.0546713e-018 ub=6.8226823e-019 uc1=-2.5583291e-010 uc=8.5033561e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094659997 voffcv=-0.16 voffl=0 vsat=84000 vth0=-0.82463101 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.066516e-008 wags=-2.0850684e-008 walpha0=-1.021993e-013 wbeta0=1.8790089e-007 wint=-1e-008 wk1=6.4792254e-008 wk2=-2.0504604e-008 wketa=-7.1778231e-009 wkt1=-1.0656933e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.6980295e-008 wtvoff=0 wu0=6.147434e-010 wua1=1.7515023e-016 wua=1.8563411e-017 wub1=-1.4365289e-025 wub=-4.6603138e-027 wuc1=3.9521569e-017 wuc=-1.2200571e-017 wvoff=-1.6325113e-009 wvth0=3.8459166e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.1 pmos a0=1.1595369 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.18927812 alpha0=7.659374e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=42.543923 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0114941 k2=-0.018959971 k3=0 k3b=0 keta=-0.0048215378 kt1=-0.3049182 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.7674521e-007 lags=1.0628082e-007 lalpha0=-3.6411844e-011 lbeta0=-5.1107814e-006 level=54 lint=0 lk1=-6.6592286e-008 lk2=-1.3552238e-009 lketa=-2.3066349e-008 lkt1=-5.8128509e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=1.230257e-007 lpdiblc2=2.5373158e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.1902635e-009 lua=8.6719409e-016 lub1=-6.1682707e-025 lub=-3.5652279e-025 luc1=-3.1520912e-017 luc=5.9904874e-017 lvoff=1.3331945e-008 lvth0=8.4932211e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.6180878e-014 pags=-2.976212e-014 palpha0=-2.3232577e-018 paramchk=1 pbeta0=8.2816979e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.26103151 pdiblc1=0.1484 pdiblc2=0.00024138051 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=2.0986491e-014 pk2=-5.9141722e-015 pketa=1.0714215e-015 pkt1=-1.5716657e-014 ppclm=-2.0904788e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-9.6149399e-017 pua=-1.6387735e-022 pub1=9.3364074e-032 pub=9.2457915e-032 puc1=3.1633858e-024 puc=-7.2547674e-024 pvag=0 pvth0=1.4780788e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010245409 ua1=1.5e-009 ua=3.5072904e-010 ub1=-2.2298632e-018 ub=1.07928e-018 uc1=-7.4455718e-011 uc=-1.5016171e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12389995 voffcv=-0.16 voffl=0 vsat=84000 vth0=-0.85684939 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=3.6902724e-008 wags=1.3597033e-008 walpha0=4.5607375e-012 wbeta0=2.5801452e-007 wint=-1e-008 wk1=-1.7315587e-008 wk2=-2.2571871e-009 wketa=-2.09262e-009 wkt1=2.3842925e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=8.0632068e-008 wtvoff=0 wu0=-2.2946106e-010 wua=-3.7369482e-017 wub1=-3.2919886e-026 wub=-1.8258434e-025 wuc1=5.7861122e-018 wuc=-6.8025157e-018 wvth0=5.5796737e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.2 pmos a0=1.2627338 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.15723172 alpha0=0.0020630943 alpha1=0 at=12000 b0=0 b1=0 beta0=44.489973 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95738704 k2=-0.012190361 k3=0 k3b=0 keta=-0.00041211629 kt1=-0.26928515 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-4.0181986e-007 lags=1.4512107e-007 lalpha0=-2.4440505e-009 lbeta0=-7.4693929e-006 level=54 lint=0 lk1=-1.0144952e-009 lk2=-9.5599917e-009 lketa=-2.8410567e-008 lkt1=-4.9000116e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.5157018e-007 lpclm=4.939508e-008 lpdiblc2=4.5176356e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.9830294e-009 lua=8.1571763e-016 lub1=3.2292957e-025 lub=-7.0271026e-026 luc1=-7.7555003e-017 luc=9.508283e-017 lvoff=-1.8520988e-008 lvoffcv=-2.2062807e-007 lvth0=-9.3166113e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9449091 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=3.2476679e-014 pags=-1.4129839e-014 palpha0=-2.2176222e-017 paramchk=1 pbeta0=-6.4121511e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32178284 pdiblc1=0.1484 pdiblc2=7.7987791e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-3.4891345e-014 pk2=8.5114085e-015 pketa=2.48312e-015 pkt1=2.4990059e-014 ppclm=7.1238421e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-6.2434711e-016 pua=-1.4935691e-022 pub1=-1.6469408e-031 pub=-3.9166112e-033 puc1=2.4194028e-023 puc=-1.7634109e-023 pvag=0 pvoff=-1.1305027e-015 pvth0=4.0552523e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0087662296 ua1=1.5e-009 ua=3.9320136e-010 ub1=-3.00524e-018 ub=8.4309868e-019 uc1=-3.6473795e-011 uc=-4.4040887e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097618657 voffcv=0.022036364 voffl=0 vsat=84000 vth0=-0.84215481 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-3.2437753e-009 wags=6.9911181e-010 walpha0=2.0941071e-011 wbeta0=3.7925089e-007 wint=-1e-008 wk1=2.8788238e-008 wk2=-1.4159481e-008 wketa=-3.2573878e-009 wkt1=-9.743475e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=4.6063177e-009 wtvoff=0 wu0=2.0634563e-010 wua=-4.9350043e-017 wub1=1.7999938e-025 wub=-1.0306741e-025 wuc1=-1.1565903e-017 wuc=1.7612973e-018 wvoff=9.3275798e-010 wvth0=3.453293e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.3 pmos a0=1.2226 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17172643 alpha0=0.0018189821 alpha1=0 at=12000 b0=0 b1=0 beta0=43.743929 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95728571 k2=-0.013145214 k3=0 k3b=0 keta=-0.0032497679 kt1=-0.27417929 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32671643 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.009064175 ua1=1.5e-009 ua=4.7467536e-010 ub1=-2.9729857e-018 ub=8.3608e-019 uc1=-4.422e-011 uc=-3.4544e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.099468536 voffcv=0 voffl=0 vsat=84000 vth0=-0.84308536 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-7.1217857e-010 walpha0=1.8726107e-011 wbeta0=3.7284643e-007 wint=-1e-008 wk1=2.5303286e-008 wk2=-1.3309361e-008 wketa=-3.0093734e-009 wkt1=-7.2474643e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=1.1721621e-008 wtvoff=0 wu0=1.4398575e-010 wua=-6.4267832e-017 wub1=1.6354971e-025 wub=-1.034586e-025 wuc1=-9.1494e-018 wvoff=8.1984321e-010 wvth0=3.8583321e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.4 pmos a0=0.68036585 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19813874 alpha0=1.233251e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=38.487806 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0017393 k2=0.015787252 k3=0 k3b=0 keta=-0.10659611 kt1=-0.33207273 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-1.1106099e-007 lags=7.4525608e-008 lalpha0=-3.2296894e-012 lbeta0=-2.9055811e-006 level=54 lint=0 lk1=-3.7831308e-008 lk2=-2.1838311e-008 lketa=2.3586916e-008 lkt1=4.5744341e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=2.9589851e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.9585121e-009 lua1=-2.7134976e-016 lua=7.9824069e-016 lub1=-3.486841e-026 lub=-3.2854766e-025 luc1=-3.6378401e-017 luc=1.3188534e-017 lvth0=-2.2948864e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-5.7518044e-014 pags=6.4820876e-015 palpha0=7.7287812e-020 paramchk=1 pbeta0=-3.6783751e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.37605618 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=1.1592273e-015 pketa=-3.6927531e-015 pkt1=-6.9014464e-015 ppclm=3.0331617e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-2.1626928e-016 pua1=1.3838838e-022 pua=-4.2295322e-023 pub1=-1.9248565e-031 pub=9.0761209e-032 puc1=3.5729363e-023 puc=-6.7906158e-024 pvag=0 pvth0=-5.4516634e-016 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0090330668 ua1=2.02998e-009 ua=-1.4390099e-010 ub1=-2.8805891e-018 ub=1.7663512e-018 uc1=7.8595636e-012 uc=8.5435958e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=84000 vth0=-0.84559037 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.969796e-007 wags=-3.0080179e-008 walpha0=-4.0713741e-013 wbeta0=1.0102328e-006 wint=-1e-008 wk2=-1.3390429e-008 wketa=1.2646415e-008 wkt1=1.4228723e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.4969243e-008 wtvoff=0 wu0=-1.4180477e-010 wua1=-2.702898e-016 wua=4.6110994e-017 wub1=2.7756517e-025 wub=-5.5754264e-025 wuc1=-9.4961592e-017 wuc=-1.2405794e-017 wvth0=1.4535189e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.5 pmos a0=1.3532832 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19095588 alpha0=0.00012387909 alpha1=0 at=12000 b0=0 b1=0 beta0=43.468326 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.977542 k2=-0.026820609 k3=0 k3b=0 keta=-0.0011314055 kt1=-0.28298126 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-4.5559467e-007 lags=7.8203234e-008 lalpha0=-6.0341539e-011 lbeta0=-5.4556076e-006 level=54 lint=0 lk1=-2.5442304e-008 lk2=-2.308677e-011 lketa=-3.0411013e-008 lkt1=-2.4677389e-008 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=-6.0780385e-008 lpdiblc2=2.5373158e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.6085514e-009 lua=5.9324665e-016 lub1=9.4139058e-026 lub=-7.4479844e-026 luc1=1.8446114e-017 luc=5.351359e-017 lvoff=1.3331945e-008 lvth0=-2.3922604e-010 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.5032345e-014 pags=-1.5442549e-014 palpha0=9.8808868e-018 paramchk=1 pbeta0=2.5867832e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.55256055 pdiblc1=0.1484 pdiblc2=0.00024138051 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-6.593562e-015 pketa=4.8172e-015 pkt1=-6.095743e-015 ppclm=7.2836314e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-3.0947618e-016 pua=-2.416415e-023 pub1=-2.6922865e-031 pub=-5.1383988e-032 puc1=-2.2319798e-023 puc=-3.9952125e-024 pvag=0 pvth0=5.9316269e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097165838 ua1=1.5e-009 ua=2.5647799e-010 ub1=-3.1325568e-018 ub=1.270125e-018 uc1=-9.9219566e-011 uc=6.6760848e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12389995 voffcv=-0.16 voffl=0 vsat=84000 vth0=-0.84960533 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-6.1907875e-008 wags=1.2741377e-008 walpha0=-1.9554792e-011 wbeta0=-2.1343096e-007 wint=-1e-008 wk2=1.7517378e-009 wketa=-3.9745875e-009 wkt1=1.2655084e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-6.8047743e-008 wtvoff=0 wu0=4.0239958e-011 wua=1.0698549e-017 wub1=4.2745384e-025 wub=-2.799153e-025 wuc1=1.8415675e-017 wuc=-1.7865566e-017 wvth0=1.8852027e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.6 pmos a0=1.1202818 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16544644 alpha0=0.0021756117 alpha1=0 at=12000 b0=0 b1=0 beta0=44.368279 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0138346 k2=-0.027555336 k3=0 k3b=0 keta=-0.0067991511 kt1=-0.33738473 kt1l=0 kt2=-0.01692062 ku0=0 kvsat=0 kvth0=0 la0=-1.7319698e-007 lags=1.0912068e-007 lalpha0=-2.5470415e-009 lbeta0=-6.5463501e-006 level=54 lint=0 lk1=-6.9428897e-008 lk2=8.6740321e-010 lketa=-2.3541705e-008 lkt1=4.1259616e-008 lkt2=4.6717994e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.5157018e-007 lpclm=2.1057807e-007 lpdiblc2=4.5176356e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.5969749e-009 lua=4.1703039e-016 lub1=-5.5513372e-025 lub=5.6792621e-026 luc1=-5.013773e-017 luc=6.0682053e-017 lvoff=-2.073766e-008 lvoffcv=-2.2062807e-007 lvth0=-1.3889719e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9449091 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-8.4120993e-014 pags=4.2303621e-015 palpha0=3.0349201e-017 paramchk=1 pbeta0=-5.3487336e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32866743 pdiblc1=0.1484 pdiblc2=7.7987791e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=3.1934371e-015 pkt1=-2.1042404e-014 pkt2=-2.3826177e-015 ppclm=-1.0964904e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=8.2540685e-017 pua=5.3973585e-023 pub1=2.831182e-031 pub=-6.8719071e-032 puc1=1.0211219e-023 puc=-8.9712851e-026 pvag=0 pvth0=1.2156213e-017 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097261353 ua1=1.5e-009 ua=4.0187094e-010 ub1=-2.5968532e-018 ub=1.1618144e-018 uc1=-4.2632236e-011 uc=7.6151064e-013 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.095789719 voffcv=0.022036364 voffl=0 vsat=84000 vth0=-0.8486567 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=6.940676e-008 wags=-3.4903977e-009 walpha0=-3.644284e-011 wbeta0=4.4131466e-007 wint=-1e-008 wk2=-6.323344e-009 wkt1=2.4987313e-008 wkt2=1.9658562e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.0951762e-009 wtvoff=0 wu0=-2.832063e-010 wua=-5.3771529e-017 wub1=-2.8277886e-026 wub=-2.6561243e-025 wuc1=-8.425098e-018 wuc=-2.1087925e-017 wvth0=6.7692544e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.7 pmos a0=1.1029829 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17634543 alpha0=0.0019212129 alpha1=0 at=12000 b0=0 b1=0 beta0=43.714429 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.0274687 k3=0 k3b=0 keta=-0.0091505 kt1=-0.33326371 kt1l=0 kt2=-0.016454 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0098856414 ua1=1.5e-009 ua=4.43524e-010 ub1=-2.6523e-018 ub=1.1674869e-018 uc1=-4.764e-011 uc=6.8224429e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=84000 vth0=-0.84879543 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=6.1004743e-008 wags=-3.0678686e-009 walpha0=-3.3411557e-011 wbeta0=3.8789143e-007 wint=-1e-008 wk2=-6.004383e-009 wkt1=2.2885594e-008 wkt2=1.72788e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wtvoff=0 wu0=-2.7496213e-010 wua=-4.838064e-017 wub=-2.724761e-025 wuc1=-7.4052e-018 wuc=-2.1096886e-017 wvth0=6.7704686e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.8 pmos a0=0.90053503 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.33423596 alpha0=9.9208915e-006 alpha1=0 at=12000 b0=0 b1=0 beta0=38.010737 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0017393 k2=0.00084217568 k3=0 k3b=0 keta=-0.090439654 kt1=-0.29527232 kt1l=0 kt2=-0.021021054 ku0=0 kvsat=0 kvth0=0 la0=-1.5725154e-007 lags=-2.5272122e-009 lalpha0=-2.4388052e-012 lbeta0=-2.5355199e-006 level=54 lint=0 lk1=-3.7831308e-008 lk2=-1.8894426e-008 lketa=1.8869231e-008 lkt1=-8.9643788e-009 lkt2=2.3228759e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=5.399252e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.9104148e-009 lua1=-1.6640984e-016 lua=6.7361745e-016 lub1=-1.373636e-025 lub=3.486153e-026 luc1=9.418752e-019 luc=-7.929225e-018 lvth0=-9.3623482e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.6274819e-015 pags=9.9716e-014 palpha0=-8.79682e-019 paramchk=1 pbeta0=-8.156116e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32055448 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-2.4028741e-015 pketa=2.0156456e-015 pkt1=4.4989585e-015 pkt2=-2.8106799e-015 ppclm=8.0438758e-016 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.5807151e-016 pua1=1.141108e-023 pua=1.0849879e-022 pub1=-6.8466478e-032 pub=-3.4896391e-031 puc1=-9.4281708e-024 puc=1.8761873e-023 pvag=0 pvth0=8.0064625e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011197346 ua1=1.8250192e-009 ua=2.9342841e-010 ub1=-2.5734555e-018 ub=9.252807e-019 uc1=-8.58396e-011 uc=1.3433638e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=84000 vth0=-0.83651091 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-6.9425106e-008 wags=-1.9475781e-007 walpha0=2.5109209e-012 wbeta0=1.5874859e-006 wint=-1e-008 wk2=4.6931134e-009 wketa=-6.902896e-009 wkt1=-3.029977e-008 wkt2=9.625616e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=8.2126294e-008 wtvoff=0 wu0=-2.7605828e-009 wua1=-2.2287265e-017 wua=-4.8305758e-016 wub1=-9.4066473e-026 wub=4.6015269e-025 wuc1=1.8414396e-017 wuc=-7.1575304e-017 wvth0=3.5490455e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.9 pmos a0=1.1841981 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20666573 alpha0=0.00011213634 alpha1=0 at=12000 b0=0 b1=0 beta0=43.288609 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.977542 k2=-0.030491622 k3=0 k3b=0 keta=-0.0062091486 kt1=-0.30256285 kt1l=0 kt2=-0.01056584 ku0=0 kvsat=0 kvth0=0 la0=-3.0248705e-007 lags=6.2788747e-008 lalpha0=-5.4773114e-011 lbeta0=-5.2377903e-006 level=54 lint=0 lk1=-2.5442304e-008 lk2=-2.8515216e-009 lketa=-2.4256788e-008 lkt1=-5.2316292e-009 lkt2=-3.0301939e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.4876612e-008 lpdiblc2=2.5373158e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.4831844e-009 lua=6.6362748e-016 lub1=-1.9632904e-025 lub=1.6080068e-026 luc1=-2.5411277e-017 luc=7.5803538e-017 lvoff=-1.8331424e-009 lvth0=-7.3771601e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.1022787e-013 pags=3.2089804e-015 palpha0=3.1430926e-018 paramchk=1 pbeta0=-4.8805786e-015 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.37742149 pdiblc1=0.1484 pdiblc2=0.00024138051 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-3.1711559e-015 pketa=-2.6294117e-015 pkt1=-2.9625112e-014 pkt2=3.6665346e-015 ppclm=-3.0808652e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.3677821e-015 pua=-1.0932496e-022 pub1=8.2237749e-032 pub=-1.6096148e-031 puc1=3.0747645e-023 puc=-3.0966051e-023 pvag=0 pvoff=1.8349755e-014 pvth0=1.4568527e-014 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010078656 ua1=1.5e-009 ua=3.1294007e-010 ub1=-2.4582886e-018 ub=9.6196324e-019 uc1=-3.43686e-011 uc=-2.9204174e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094280644 voffcv=-0.16 voffl=0 vsat=84000 vth0=-0.84038823 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.4268502e-007 wags=-6.2675398e-009 walpha0=-5.3460607e-012 wbeta0=4.02688e-009 wint=-1e-008 wk2=6.1936639e-009 wketa=2.1694816e-009 wkt1=3.6348805e-008 wkt2=-3.0251936e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.4387051e-007 wtvoff=0 wu0=-3.9786675e-010 wua=-5.7620563e-017 wub1=-3.8841067e-025 wub=9.2960446e-026 wuc1=-6.0053994e-017 wuc=2.5549547e-017 wvoff=-3.5839366e-008 wvth0=-9.2674868e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.10 pmos a0=1.1835318 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16674407 alpha0=0.0021451803 alpha1=0 at=12000 b0=0 b1=0 beta0=44.168746 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0138346 k2=-0.036023613 k3=0 k3b=0 keta=-0.0067991511 kt1=-0.29671705 kt1l=0 kt2=-0.012759382 ku0=0 kvsat=0 kvth0=0 la0=-3.0167941e-007 lags=1.111738e-007 lalpha0=-2.5188225e-009 lbeta0=-6.3045161e-006 level=54 lint=0 lk1=-6.9428897e-008 lk2=3.853252e-009 lketa=-2.3541705e-008 lkt1=-1.2316734e-008 lkt2=-3.7162041e-010 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.5157018e-007 lpclm=6.6528672e-008 lpdiblc2=4.5176356e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.3317214e-009 lua1=1.2610963e-016 lua=2.3441974e-016 lub1=4.4158364e-026 luc1=1.3638952e-017 luc=6.0607911e-017 lvoff=2.8514282e-009 lvoffcv=-2.2062807e-007 lvth0=-4.5159809e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9449091 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.1342757e-014 pags=1.746085e-015 palpha0=-3.795837e-018 paramchk=1 pbeta0=-8.2749248e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34305511 pdiblc1=0.1484 pdiblc2=7.7987791e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-4.1943999e-016 pkt1=4.378498e-014 pkt2=3.7199203e-015 ppclm=1.6333487e-013 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=4.0349748e-016 pua1=-1.5259265e-022 pua=2.7493248e-022 pub1=-4.4202522e-031 puc1=-6.6958565e-023 pvag=0 pvoff=-2.8542797e-014 pvth0=3.795837e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011028707 ua1=1.3959491e-009 ua=6.6707187e-010 ub1=-2.6567105e-018 ub=9.7523062e-019 uc1=-6.658826e-011 uc=-1.6666527e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.098145801 voffcv=0.022036364 voffl=0 vsat=84000 vth0=-0.84274894 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-7.1257249e-009 wags=-5.0605305e-009 walpha0=3.7912875e-013 wbeta0=6.8274957e-007 wint=-1e-008 wk2=3.9232712e-009 wkt1=-2.4220578e-008 wkt2=-3.0692412e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=-1.631391e-008 wtvoff=0 wu0=-1.8593186e-009 wua1=1.2590153e-016 wua=-3.7466465e-016 wub1=4.4149543e-026 wub=-3.9846056e-026 wuc1=2.0561691e-017 wvoff=2.8508586e-009 wvth0=-3.7912875e-010 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.11 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17784813 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.53905 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.03563875 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29794725 kt1l=0 kt2=-0.0127965 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.01116172 ua1=1.408545e-009 ua=6.9048575e-010 ub1=-2.6523e-018 ub=9.7523062e-019 uc1=-6.5226e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=84000 vth0=-0.8432 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-4.8861312e-009 wbeta0=6.000995e-007 wint=-1e-008 wk2=3.8813775e-009 wkt1=-1.9847327e-008 wkt2=-2.697695e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wtvoff=0 wu0=-1.8190172e-009 wua1=1.1066055e-016 wua=-3.4720436e-016 wub=-3.9846056e-026 wuc1=1.387386e-017 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.12 pmos a0=0.89359946 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.31477964 alpha0=1.0171733e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=38.169327 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0017393 k2=0.0013110182 k3=0 k3b=0 keta=-0.091129254 kt1=-0.29829927 kt1l=0 kt2=-0.020059454 ku0=0 kvsat=0 kvth0=0 la0=-1.5741412e-007 lags=7.4344262e-009 lalpha0=-2.5266856e-012 lbeta0=-2.6169996e-006 level=54 lint=0 lk1=-3.7831308e-008 lk2=-1.9134473e-008 lketa=1.9070594e-008 lkt1=-8.5149324e-009 lkt2=2.0420887e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=5.4072878e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.8946234e-009 lua1=-1.6526988e-016 lua=6.844565e-016 lub1=-1.442034e-025 luc=-6.054912e-018 lvth0=-8.5625018e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32875891 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010921564 ua1=1.8227927e-009 ua=2.4517091e-010 ub1=-2.5828527e-018 ub=9.7125e-019 uc1=-8.4e-011 uc=1.27186e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=84000 vth0=-0.83615636 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.13 pmos a0=1.1984524 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.2060396 alpha0=0.00011160227 alpha1=0 at=12000 b0=0 b1=0 beta0=43.289011 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.977542 k2=-0.029872874 k3=0 k3b=0 keta=-0.0059924171 kt1=-0.2989316 kt1l=0 kt2=-0.010868057 ku0=0 kvsat=0 kvth0=0 la0=-3.1349883e-007 lags=6.3109325e-008 lalpha0=-5.4459119e-011 lbeta0=-5.2382779e-006 level=54 lint=0 lk1=-2.5442304e-008 lk2=-3.1683204e-009 lketa=-2.4519466e-008 lkt1=-8.1911808e-009 lkt2=-2.6639067e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.1798824e-008 lpdiblc2=2.5373158e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.3465428e-009 lua=6.5270591e-016 lub1=-1.8811348e-025 luc1=-2.2339584e-017 luc=7.2710027e-017 lvth0=-5.9217627e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.39179417 pdiblc1=0.1484 pdiblc2=0.00024138051 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010038909 ua1=1.5e-009 ua=3.0718377e-010 ub1=-2.4970909e-018 ub=9.7125e-019 uc1=-4.0368e-011 uc=-2.6651771e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=84000 vth0=-0.84131406 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.14 pmos a0=1.1828199 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16623852 alpha0=0.0021452182 alpha1=0 at=12000 b0=0 b1=0 beta0=44.236953 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0138346 k2=-0.035631678 k3=0 k3b=0 keta=-0.0067991511 kt1=-0.29913669 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.9455227e-007 lags=1.1134823e-007 lalpha0=-2.5192017e-009 lbeta0=-6.3871827e-006 level=54 lint=0 lk1=-6.9428897e-008 lk2=3.81135e-009 lketa=-2.3541705e-008 lkt1=-7.9426106e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.5157018e-007 lpclm=8.2845841e-008 lpdiblc2=4.5176356e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.3720308e-009 lua1=1.1086561e-016 lua=2.6188552e-016 luc1=6.9497843e-018 luc=6.0607911e-017 lvoffcv=-2.2062807e-007 lvth0=-4.1367764e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9449091 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34142534 pdiblc1=0.1484 pdiblc2=7.7987791e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010842961 ua1=1.4085267e-009 ua=6.2964284e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.4534145e-011 uc=-1.6666527e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0.022036364 voffl=0 vsat=84000 vth0=-0.84278682 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.model pmos_3p3.15 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17736 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.599 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.4e-011 cgdo=1.364e-010 cgidl=7.5 cgsl=4.4e-011 cgso=1.364e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035251 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29993 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.3e-009 toxm=7.9e-009 toxp=8.3e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.01098 ua1=1.4196e-009 ua=6.558e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.384e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=84000 vth0=-0.8432 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=1.2e-008 xpart=0 xtis=3 xw=-1e-008
.subckt pplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 par=1 r_rsh0='rsh_pplus_u_m' r_dw=2.75e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.375e-3 r_tc2=1e-6 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model pn_junction d cj=0.00094344 level=2
d1 1 3 pn_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends pplus_u_m1
.endl pmos_3p3_s

.lib pmos_3p3_fs
.subckt pmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.00666
.param par_k=0.002833
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b pplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b pplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b pmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model pmos_3p3.0 pmos a0=1.039392 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.18391438 alpha0=1.1653153e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=39.988812 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.87205009 k2=0.029903393 k3=0 k3b=0 keta=-0.067178738 kt1=-0.28327726 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.1366429e-007 lags=1.0913958e-007 lalpha0=-3.1380589e-012 lbeta0=-3.7819465e-006 level=54 lint=0 lk1=4.25291e-009 lk2=-2.5868222e-008 lketa=8.7913147e-009 lkt1=-1.6612629e-008 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=7.4286569e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.5375194e-009 lua1=1.7581418e-016 lua=1.0774293e-015 lub1=-6.9766226e-025 lub=-1.5002929e-025 luc1=6.0619732e-017 luc=8.6809692e-018 lvoff=-1.6386998e-009 lvth0=-7.9299856e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.7738176e-015 pags=-1.2242165e-014 palpha0=6.4786605e-020 paramchk=1 pbeta0=1.1986341e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.35338606 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-2.1256353e-014 pk2=3.4616668e-015 pketa=3.7105918e-015 pkt1=1.9661049e-015 ppclm=6.6284179e-015 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-5.3349279e-016 pua1=-9.0544304e-023 pua=-1.9437706e-022 pub1=1.515108e-031 pub=1.3739739e-033 puc1=-1.4245637e-023 puc=-4.5344012e-024 pvag=0 pvoff=8.439304e-016 pvth0=2.388645e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0075928117 ua1=1.1539091e-009 ua=-6.122012e-011 ub1=-2.0676223e-018 ub=6.7836503e-019 uc1=-2.5586018e-010 uc=8.579096e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094635213 voffcv=-0.16 voffl=0 vsat=90000 vth0=-0.81501176 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.0928007e-008 wags=-2.1847527e-008 walpha0=-1.0367347e-013 wbeta0=1.9714501e-007 wint=-1e-008 wk1=6.6268653e-008 wk2=-2.1061108e-008 wketa=-7.3043146e-009 wkt1=-1.0941603e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.8018309e-008 wtvoff=0 wu0=6.1967943e-010 wua1=1.7823682e-016 wua=1.383858e-017 wub1=-1.440724e-025 wub=-4.7707426e-027 wuc1=4.0387143e-017 wuc=-1.2711987e-017 wvoff=-1.6612803e-009 wvth0=4.0333546e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.1 pmos a0=1.1561845 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.1893918 alpha0=7.6165264e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=42.499959 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0117972 k2=-0.018870868 k3=0 k3b=0 keta=-0.0048813173 kt1=-0.30596768 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.7299485e-007 lags=1.0635705e-007 lalpha0=-3.5910211e-011 lbeta0=-5.0576089e-006 level=54 lint=0 lk1=-6.6738621e-008 lk2=-1.0908973e-009 lketa=-2.2855775e-008 lkt1=-5.0858969e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=1.2254291e-007 lpdiblc2=2.5091844e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.18112e-009 lua=8.6448742e-016 lub1=-6.1392387e-025 lub=-3.564674e-025 luc1=-3.1304785e-017 luc=5.9546517e-017 lvoff=1.3184133e-008 lvth0=8.3367507e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.6509626e-014 pags=-3.0366798e-014 palpha0=-2.3704594e-018 paramchk=1 pbeta0=8.4499576e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.25839327 pdiblc1=0.1484 pdiblc2=0.00024301606 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=2.1412875e-014 pk2=-6.0343307e-015 pketa=1.0931896e-015 pkt1=-1.6035973e-014 ppclm=-2.1329512e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-9.8102871e-017 pua=-1.6720685e-022 pub1=9.5260957e-032 pub=9.4336388e-032 puc1=3.2276564e-024 puc=-7.4021628e-024 pvag=0 pvth0=1.508109e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010262889 ua1=1.5e-009 ua=3.5795686e-010 ub1=-2.2324617e-018 ub=1.0847393e-018 uc1=-7.4906407e-011 uc=-1.4338071e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12381402 voffcv=-0.16 voffl=0 vsat=90000 vth0=-0.84703289 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=3.7967e-008 wags=1.3830885e-008 walpha0=4.6901179e-012 wbeta0=2.6675886e-007 wint=-1e-008 wk1=-1.772589e-008 wk2=-2.3681999e-009 wketa=-2.151948e-009 wkt1=2.4495559e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=8.3053604e-008 wtvoff=0 wu0=-2.3738733e-010 wua=-3.9646086e-017 wub1=-3.3344363e-026 wub=-1.8776762e-025 wuc1=5.9908956e-018 wuc=-7.0667866e-018 wvth0=5.7666931e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.2 pmos a0=1.2627392 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.15724995 alpha0=0.0020613963 alpha1=0 at=12000 b0=0 b1=0 beta0=44.471345 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95616008 k2=-0.011590073 k3=0 k3b=0 keta=-0.00028266778 kt1=-0.26888633 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-4.0171294e-007 lags=1.451844e-007 lalpha0=-2.4340693e-009 lbeta0=-7.439044e-006 level=54 lint=0 lk1=4.7102587e-010 lk2=-9.886097e-009 lketa=-2.8410943e-008 lkt1=-4.9880168e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4953018e-007 lpclm=4.6187031e-008 lpdiblc2=4.500927e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.9985114e-009 lua=8.1904358e-016 lub1=3.2872945e-025 lub=-6.9844795e-026 luc1=-7.8295637e-017 luc=9.548005e-017 lvoff=-1.8404477e-008 lvoffcv=-2.1981207e-007 lvth0=-9.4543724e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9450909 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=3.3384084e-014 pags=-1.452463e-014 palpha0=-2.279583e-017 paramchk=1 pbeta0=-6.5913079e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32160177 pdiblc1=0.1484 pdiblc2=7.8136709e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-3.5866216e-014 pk2=8.7492189e-015 pketa=2.5524988e-015 pkt1=2.5688286e-014 ppclm=7.3228837e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-6.4179149e-016 pua=-1.5352997e-022 pub1=-1.6929566e-031 pub=-4.0260421e-033 puc1=2.4870014e-023 puc=-1.8126809e-023 pvag=0 pvoff=-1.1620891e-015 pvth0=4.1685569e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0087584261 ua1=1.5e-009 ua=3.9557594e-010 ub1=-3.0128038e-018 ub=8.474689e-019 uc1=-3.6006695e-011 uc=-4.4084373e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097664506 voffcv=0.021963636 voffl=0 vsat=90000 vth0=-0.83230514 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-3.3357398e-009 wags=7.1650729e-010 walpha0=2.1598538e-011 wbeta0=3.9127265e-007 wint=-1e-008 wk1=2.9690576e-008 wk2=-1.4606238e-008 wketa=-3.3599854e-009 wkt1=-1.0044391e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=4.7768253e-009 wtvoff=0 wu0=2.1268603e-010 wua=-5.0968009e-017 wub1=1.8565946e-025 wub=-1.0634177e-025 wuc1=-1.1924963e-017 wuc=1.8112319e-018 wvoff=9.6199433e-010 wvth0=3.5643356e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.3 pmos a0=1.2226 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17175679 alpha0=0.0018181839 alpha1=0 at=12000 b0=0 b1=0 beta0=43.728036 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95620714 k2=-0.012577893 k3=0 k3b=0 keta=-0.0031214911 kt1=-0.27387036 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32621679 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0090580375 ua1=1.5e-009 ua=4.7741482e-010 ub1=-2.9799571e-018 ub=8.4049e-019 uc1=-4.383e-011 uc=-3.4544e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.099503482 voffcv=0 voffl=0 vsat=90000 vth0=-0.83324982 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-7.3479464e-010 walpha0=1.9320777e-011 wbeta0=3.8468661e-007 wint=-1e-008 wk1=2.6106821e-008 wk2=-1.3732015e-008 wketa=-3.1049396e-009 wkt1=-7.4776161e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=1.2093855e-008 wtvoff=0 wu0=1.4855819e-010 wua=-6.6308733e-017 wub1=1.6874343e-025 wub=-1.0674405e-025 wuc1=-9.43995e-018 wvoff=8.458783e-010 wvth0=3.980858e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.4 pmos a0=0.67581086 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.200375 alpha0=1.2249381e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=38.401961 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0007271 k2=0.015311208 k3=0 k3b=0 keta=-0.1060667 kt1=-0.33217428 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-1.0822777e-007 lags=7.2879057e-008 lalpha0=-3.1611736e-012 lbeta0=-2.8404732e-006 level=54 lint=0 lk1=-3.7021562e-008 lk2=-2.1380073e-008 lketa=2.3111339e-008 lkt1=5.0237373e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=2.8716008e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.9183067e-009 lua1=-2.6663904e-016 lua=7.8149042e-016 lub1=-3.2595866e-026 lub=-3.2223504e-025 luc1=-3.5883051e-017 luc=1.2960088e-017 lvth0=-2.2414438e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-5.7073625e-014 pags=6.4320031e-015 palpha0=7.669064e-020 paramchk=1 pbeta0=-3.6499537e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.37672 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=1.1502704e-015 pketa=-3.6642206e-015 pkt1=-6.8481216e-015 ppclm=3.0097257e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-2.1459826e-016 pua1=1.3731911e-022 pua=-4.1968523e-023 pub1=-1.9099839e-031 pub=9.0059933e-032 puc1=3.5453296e-023 puc=-6.7381475e-024 pvag=0 pvth0=-5.4095405e-016 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0090866629 ua1=2.02488e-009 ua=-1.2290839e-010 ub1=-2.8837292e-018 ub=1.7620586e-018 uc1=7.6479273e-012 uc=8.5890808e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=90000 vth0=-0.83576942 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.9817231e-007 wags=-3.0324746e-008 walpha0=-4.1073109e-013 wbeta0=1.0143734e-006 wint=-1e-008 wk2=-1.3546134e-008 wketa=1.2722988e-008 wkt1=1.4240363e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.6001332e-008 wtvoff=0 wu0=-1.4965392e-010 wua1=-2.703132e-016 wua=4.5608039e-017 wub1=2.7622264e-025 wub=-5.6287295e-025 wuc1=-9.5319534e-017 wuc=-1.2763408e-017 wvth0=1.4723553e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.5 pmos a0=1.3508441 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19135754 alpha0=0.00012364806 alpha1=0 at=12000 b0=0 b1=0 beta0=43.434876 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.977378 k2=-0.026834606 k3=0 k3b=0 keta=-0.0012954815 kt1=-0.28324255 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-4.5114467e-007 lags=7.7459926e-008 lalpha0=-5.9751701e-011 lbeta0=-5.3971937e-006 level=54 lint=0 lk1=-2.5160224e-008 lk2=3.0000655e-011 lketa=-3.0112442e-008 lkt1=-2.4354946e-008 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=-6.0690117e-008 lpdiblc2=2.5091844e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.593197e-009 lua=5.8686291e-016 lub1=9.525255e-026 lub=-7.3242364e-026 luc1=1.842044e-017 luc=5.2952294e-017 lvoff=1.3184133e-008 lvth0=-2.8410138e-010 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.5237532e-014 pags=-1.5484779e-014 palpha0=9.9079077e-018 paramchk=1 pbeta0=2.5938572e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.55271631 pdiblc1=0.1484 pdiblc2=0.00024301606 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-6.6115932e-015 pketa=4.8303734e-015 pkt1=-6.1124128e-015 ppclm=7.3035497e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-3.103225e-016 pua=-2.4230231e-023 pub1=-2.699649e-031 pub=-5.1524505e-032 puc1=-2.2380835e-023 puc=-4.006138e-024 pvag=0 pvth0=5.9478478e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097266426 ua1=1.5e-009 ua=2.6021662e-010 ub1=-3.1353993e-018 ub=1.2719156e-018 uc1=-9.9248709e-011 uc=7.1659939e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12381402 voffcv=-0.16 voffl=0 vsat=90000 vth0=-0.83962246 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-6.2282725e-008 wags=1.2818526e-008 walpha0=-1.9763521e-011 wbeta0=-2.1472328e-007 wint=-1e-008 wk2=1.7331254e-009 wketa=-3.9986535e-009 wkt1=1.2792118e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-6.8522762e-008 wtvoff=0 wu0=3.8779626e-011 wua=1.0690141e-017 wub1=4.3166852e-025 wub=-2.8416343e-025 wuc1=1.8527181e-017 wuc=-1.814138e-017 wvth0=1.950321e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.6 pmos a0=1.1196626 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16551068 alpha0=0.0021750673 alpha1=0 at=12000 b0=0 b1=0 beta0=44.362547 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0138117 k2=-0.027503825 k3=0 k3b=0 keta=-0.0068069114 kt1=-0.33757353 kt1l=0 kt2=-0.016935002 ku0=0 kvsat=0 kvth0=0 la0=-1.7187734e-007 lags=1.0868294e-007 lalpha0=-2.5378662e-009 lbeta0=-6.5178205e-006 level=54 lint=0 lk1=-6.9172112e-008 lk2=8.3841624e-010 lketa=-2.3454635e-008 lkt1=4.127688e-008 lkt2=4.6737542e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4953018e-007 lpclm=2.0988775e-007 lpdiblc2=4.500927e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.5904022e-009 lua=4.150523e-016 lub1=-5.55366e-025 lub=5.7137303e-026 luc1=-5.0034723e-017 luc=6.0458343e-017 lvoff=-2.0660961e-008 lvoffcv=-2.1981207e-007 lvth0=-1.3839329e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9450909 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-8.4981251e-014 pags=4.2736236e-015 palpha0=3.0659565e-017 paramchk=1 pbeta0=-5.4034322e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.328728 pdiblc1=0.1484 pdiblc2=7.8136709e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=3.2260946e-015 pkt1=-2.1257593e-014 pkt2=-2.4069834e-015 ppclm=-1.1077036e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=8.3384782e-017 pua=5.4525543e-023 pub1=2.8601349e-031 pub=-6.9421823e-032 puc1=1.0315643e-023 puc=-9.0630294e-026 pvag=0 pvth0=1.2280528e-017 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097289562 ua1=1.5e-009 ua=4.0244395e-010 ub1=-2.5968078e-018 ub=1.1639854e-018 uc1=-4.2580527e-011 uc=9.5237707e-013 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.095796556 voffcv=0.021963636 voffl=0 vsat=90000 vth0=-0.838712 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=7.0348718e-008 wags=-3.5377679e-009 walpha0=-3.6942045e-011 wbeta0=4.4730399e-007 wint=-1e-008 wk2=-6.4106558e-009 wkt1=2.5329519e-008 wkt2=1.9925359e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.1068181e-009 wtvoff=0 wu0=-2.8713699e-010 wua=-5.4505036e-017 wub1=-2.8578486e-026 wub=-2.6934777e-025 wuc1=-8.5394397e-018 wuc=-2.1382694e-017 wvth0=6.8638701e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.7 pmos a0=1.1024886 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17637029 alpha0=0.0019214836 alpha1=0 at=12000 b0=0 b1=0 beta0=43.711286 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.02742005 k3=0 k3b=0 keta=-0.0091505 kt1=-0.33344914 kt1l=0 kt2=-0.016468 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0098878693 ua1=1.5e-009 ua=4.43916e-010 ub1=-2.6523e-018 ub=1.1696946e-018 uc1=-4.758e-011 uc=6.9933786e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=90000 vth0=-0.83885029 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=6.1857386e-008 wags=-3.1107471e-009 walpha0=-3.3878539e-011 wbeta0=3.9331286e-007 wint=-1e-008 wk2=-6.0883043e-009 wkt1=2.3205459e-008 wkt2=1.75203e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wtvoff=0 wu0=-2.7880518e-010 wua=-4.905684e-017 wub=-2.762844e-025 wuc1=-7.5087e-018 wuc=-2.139175e-017 wvth0=6.8650971e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.8 pmos a0=0.89635642 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.33424764 alpha0=9.8546141e-006 alpha1=0 at=12000 b0=0 b1=0 beta0=37.942253 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0007271 k2=0.0003347419 k3=0 k3b=0 keta=-0.089931978 kt1=-0.29549971 kt1l=0 kt2=-0.020962848 ku0=0 kvsat=0 kvth0=0 la0=-1.5388505e-007 lags=-2.5134022e-009 lalpha0=-2.3862494e-012 lbeta0=-2.4809199e-006 level=54 lint=0 lk1=-3.7021562e-008 lk2=-1.8489037e-008 lketa=1.8464538e-008 lkt1=-8.7743217e-009 lkt2=2.2742923e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=5.2836533e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.8695879e-009 lua1=-1.628526e-016 lua=6.5915544e-016 lub1=-1.3439579e-025 lub=3.4256322e-026 luc1=9.2552394e-019 luc=-7.7670863e-018 lvth0=-9.1651899e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.6000271e-015 pags=9.8033842e-014 palpha0=-8.6484221e-019 paramchk=1 pbeta0=-8.0185264e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32196515 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-2.3623388e-015 pketa=1.9816427e-015 pkt1=4.4230633e-015 pkt2=-2.7632651e-015 ppclm=7.9081797e-016 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.5540493e-016 pua1=1.121858e-023 pua=1.0666847e-022 pub1=-6.7311483e-032 pub=-3.4307707e-031 puc1=-9.2691223e-024 puc=1.8445369e-023 pvag=0 pvth0=7.8713975e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011249601 ua1=1.820576e-009 ua=3.1164935e-010 ub1=-2.5770911e-018 ub=9.2602732e-019 uc1=-8.5821897e-011 uc=1.3415357e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=90000 vth0=-0.82676296 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-6.9790553e-008 wags=-1.9298e-007 walpha0=2.4989109e-012 wbeta0=1.5729191e-006 wint=-1e-008 wk2=4.6502732e-009 wketa=-6.8807038e-009 wkt1=-3.0319244e-008 wkt2=9.5946705e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=8.2528472e-008 wtvoff=0 wu0=-2.7776236e-009 wua1=-2.208382e-017 wua=-4.8237961e-016 wub1=-9.6342676e-026 wub=4.5290511e-025 wuc1=1.8246304e-017 wuc=-7.1402667e-017 wvth0=3.7806977e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.9 pmos a0=1.1821897 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20707304 alpha0=0.00011178547 alpha1=0 at=12000 b0=0 b1=0 beta0=43.254845 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.977378 k2=-0.030512551 k3=0 k3b=0 keta=-0.0063663954 kt1=-0.3026115 kt1l=0 kt2=-0.010584133 ku0=0 kvsat=0 kvth0=0 la0=-2.9908837e-007 lags=6.2091296e-008 lalpha0=-5.4167125e-011 lbeta0=-5.1797167e-006 level=54 lint=0 lk1=-2.5160224e-008 lk2=-2.818612e-009 lketa=-2.3986778e-008 lkt1=-5.1615319e-009 lkt2=-2.9980948e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.4613381e-008 lpdiblc2=2.5091844e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.4562116e-009 lua=6.5631445e-016 lub1=-1.941859e-025 lub=1.5967497e-026 luc1=-2.5142093e-017 luc=7.4975743e-017 lvoff=-1.8203092e-009 lvth0=-7.3013165e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.0951088e-013 pags=3.1881072e-015 palpha0=3.122648e-018 paramchk=1 pbeta0=-4.8488322e-015 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.37752254 pdiblc1=0.1484 pdiblc2=0.00024301606 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-3.1505287e-015 pketa=-2.6123084e-015 pkt1=-2.9432412e-014 pkt2=3.6426852e-015 ppclm=-3.0608253e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.3588852e-015 pua=-1.0861384e-022 pub1=8.1702823e-032 pub=-1.5991449e-031 puc1=3.0547643e-023 puc=-3.0764628e-023 pvag=0 pvoff=1.8230397e-014 pvth0=1.4473764e-014 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.01009483 ua1=1.5e-009 ua=3.1724186e-010 ub1=-2.459394e-018 ub=9.6202895e-019 uc1=-3.4507691e-011 uc=-2.8726012e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094277714 voffcv=-0.16 voffl=0 vsat=90000 vth0=-0.830432 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.4263238e-007 wags=-6.2758015e-009 walpha0=-5.3504792e-012 wbeta0=4.013934e-009 wint=-1e-008 wk2=6.2018282e-009 wketa=2.1625069e-009 wkt1=3.6325391e-008 wkt2=-3.0154679e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.4433767e-007 wtvoff=0 wu0=-4.0856791e-010 wua=-5.8595534e-017 wub1=-3.8967792e-025 wub=9.2348847e-026 wuc1=-6.0133156e-017 wuc=2.5467408e-017 wvoff=-3.5886608e-008 wvth0=-9.2160872e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.10 pmos a0=1.1834353 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16678281 alpha0=0.0021443499 alpha1=0 at=12000 b0=0 b1=0 beta0=44.166386 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0138117 k2=-0.036023963 k3=0 k3b=0 keta=-0.0068069114 kt1=-0.29671112 kt1l=0 kt2=-0.012758239 ku0=0 kvsat=0 kvth0=0 la0=-3.0059299e-007 lags=1.107619e-007 lalpha0=-2.509505e-009 lbeta0=-6.2808583e-006 level=54 lint=0 lk1=-6.9172112e-008 lk2=3.8391732e-009 lketa=-2.3454635e-008 lkt1=-1.2289189e-008 lkt2=-3.717759e-010 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4953018e-007 lpclm=6.6215436e-008 lpdiblc2=4.500927e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.32663e-009 lua1=1.2570597e-016 lua=2.3343966e-016 lub1=4.4176841e-026 luc1=1.3616046e-017 luc=6.038375e-017 lvoff=2.8526213e-009 lvoffcv=-2.1981207e-007 lvth0=-4.5008395e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9450909 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.1408259e-014 pags=1.7476882e-015 palpha0=-3.7993221e-018 paramchk=1 pbeta0=-8.2825222e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34308375 pdiblc1=0.1484 pdiblc2=7.8136709e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-4.1982509e-016 pkt1=4.382518e-014 pkt2=3.7233357e-015 ppclm=1.6348483e-013 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=4.0386794e-016 pua1=-1.5273275e-022 pua=2.751849e-022 pub1=-4.4243106e-031 puc1=-6.7020042e-023 pvag=0 pvoff=-2.8569002e-014 pvth0=3.7993221e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011029914 ua1=1.3959388e-009 ua=6.6730377e-010 ub1=-2.6567142e-018 ub=9.7524707e-019 uc1=-6.6592244e-011 uc=-1.6646548e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.098146034 voffcv=0.021963636 voffl=0 vsat=90000 vth0=-0.83275028 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-7.1351178e-009 wags=-5.0834017e-009 walpha0=3.7962851e-013 wbeta0=6.8563925e-007 wint=-1e-008 wk2=3.941312e-009 wkt1=-2.4318311e-008 wkt2=-3.0822315e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=-1.6335415e-008 wtvoff=0 wu0=-1.8678007e-009 wua1=1.2643439e-016 wua=-3.7630972e-016 wub1=4.420774e-026 wub=-4.0030695e-026 wuc1=2.0634796e-017 wvoff=2.8546166e-009 wvth0=-3.7962851e-010 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.11 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17785014 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.538802 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035640352 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29793906 kt1l=0 kt2=-0.012795386 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011162471 ua1=1.4084993e-009 ua=6.9062908e-010 ub1=-2.6523e-018 ub=9.7524707e-019 uc1=-6.5231727e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=90000 vth0=-0.8332 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-4.9087726e-009 wbeta0=6.0288024e-007 wint=-1e-008 wk2=3.899363e-009 wkt1=-1.9939296e-008 wkt2=-2.7101956e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wtvoff=0 wu0=-1.8274461e-009 wua1=1.1117333e-016 wua=-3.4881323e-016 wub=-4.0030695e-026 wuc1=1.3938149e-017 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.12 pmos a0=0.88938782 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.31497855 alpha0=1.0104131e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=38.099309 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0007271 k2=0.00079907273 k3=0 k3b=0 keta=-0.090619018 kt1=-0.29852709 kt1l=0 kt2=-0.020004818 ku0=0 kvsat=0 kvth0=0 la0=-1.5404481e-007 lags=7.2752989e-009 lalpha0=-2.4726041e-012 lbeta0=-2.560985e-006 level=54 lint=0 lk1=-3.7021562e-008 lk2=-1.8724917e-008 lketa=1.8662405e-008 lkt1=-8.3326778e-009 lkt2=1.9983796e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=5.2915497e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.8540707e-009 lua1=-1.6173242e-016 lua=6.6980631e-016 lub1=-1.4111686e-025 luc=-5.925312e-018 lvth0=-8.3792291e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.33020564 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010972255 ua1=1.8183709e-009 ua=2.6348364e-010 ub1=-2.5867109e-018 ub=9.7125e-019 uc1=-8.4e-011 uc=1.27024e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=90000 vth0=-0.82638545 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.13 pmos a0=1.1964316 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.2064464 alpha0=0.00011125123 alpha1=0 at=12000 b0=0 b1=0 beta0=43.255246 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.977378 k2=-0.029893297 k3=0 k3b=0 keta=-0.0061504686 kt1=-0.2989844 kt1l=0 kt2=-0.010885229 ku0=0 kvsat=0 kvth0=0 la0=-3.1002305e-007 lags=6.2409629e-008 lalpha0=-5.3855328e-011 lbeta0=-5.1802008e-006 level=54 lint=0 lk1=-2.5160224e-008 lk2=-3.133193e-009 lketa=-2.4247618e-008 lkt1=-8.1003648e-009 lkt2=-2.6343719e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.155714e-008 lpdiblc2=2.5091844e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.3205266e-009 lua=6.4546933e-016 lub1=-1.8602786e-025 luc1=-2.2091904e-017 luc=7.1903887e-017 lvth0=-5.8561079e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.39193469 pdiblc1=0.1484 pdiblc2=0.00024301606 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010054034 ua1=1.5e-009 ua=3.1139109e-010 ub1=-2.4983034e-018 ub=9.7125e-019 uc1=-4.0512e-011 uc=-2.6183086e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=90000 vth0=-0.83135223 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.14 pmos a0=1.1827228 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16627523 alpha0=0.0021443878 alpha1=0 at=12000 b0=0 b1=0 beta0=44.234847 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0138117 k2=-0.035630422 k3=0 k3b=0 keta=-0.0068069114 kt1=-0.29913931 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.9346286e-007 lags=1.109364e-007 lalpha0=-2.5098843e-009 lbeta0=-6.3635595e-006 level=54 lint=0 lk1=-6.9172112e-008 lk2=3.7972536e-009 lketa=-2.3454635e-008 lkt1=-7.9132346e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4953018e-007 lpclm=8.2539433e-008 lpdiblc2=4.500927e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.3669563e-009 lua1=1.1045557e-016 lua=2.6091693e-016 luc1=6.9240803e-018 luc=6.038375e-017 lvoffcv=-2.1981207e-007 lvth0=-4.1214764e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9450909 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34145265 pdiblc1=0.1484 pdiblc2=7.8136709e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010843414 ua1=1.4085633e-009 ua=6.2972916e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.4531855e-011 uc=-1.6646548e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0.021963636 voffl=0 vsat=90000 vth0=-0.83278818 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.model pmos_3p3.15 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17736 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.599 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4.2e-011 cgdo=1.302e-010 cgidl=7.5 cgsl=4.2e-011 cgso=1.302e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035251 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29993 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=8.1e-009 toxm=7.9e-009 toxp=8.1e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.01098 ua1=1.4196e-009 ua=6.558e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.384e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=90000 vth0=-0.8332 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=8e-009 xpart=0 xtis=3 xw=-5e-009
.subckt pplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 par=1 r_rsh0='rsh_pplus_u_m' r_dw=2.75e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.375e-3 r_tc2=1e-6 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model pn_junction d cj=0.00094344 level=2
d1 1 3 pn_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends pplus_u_m1
.endl pmos_3p3_fs

.lib pmos_3p3_sf
.subckt pmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.00666
.param par_k=0.002833
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b pplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b pplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b pmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model pmos_3p3.0 pmos a0=1.0151475 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19776586 alpha0=1.1317951e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=39.557841 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.86723166 k2=0.028783357 k3=0 k3b=0 keta=-0.0656473 kt1=-0.28420773 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-1.9522869e-007 lags=1.0075502e-007 lalpha0=-2.8752733e-012 lbeta0=-3.4683987e-006 level=54 lint=0 lk1=5.4966687e-009 lk2=-2.3923245e-008 lketa=7.7609556e-009 lkt1=-1.5344138e-008 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=6.7448817e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.3613853e-009 lua1=1.6766018e-016 lua=1.0002135e-015 lub1=-6.4960147e-025 lub=-1.3733536e-025 luc1=5.6525433e-017 luc=8.2831734e-018 lvoff=-1.5626994e-009 lvth0=-7.4340753e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.6965346e-015 pags=-1.1901079e-014 palpha0=6.2981547e-020 paramchk=1 pbeta0=1.1652383e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.35913516 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-2.0664117e-014 pk2=3.3652193e-015 pketa=3.6072088e-015 pkt1=1.9113261e-015 ppclm=6.4437396e-015 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-5.1862883e-016 pua1=-8.8021596e-023 pua=-1.8896141e-022 pub1=1.4728947e-031 pub=1.3356928e-033 puc1=-1.3848731e-023 puc=-4.4080656e-024 pvag=0 pvoff=8.2041716e-016 pvth0=2.3220935e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0078239364 ua1=1.1592273e-009 ua=5.7221977e-011 ub1=-2.1333843e-018 ub=6.6233941e-019 uc1=-2.5243909e-010 uc=8.7831657e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094684782 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.68623384 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.1291855e-008 wags=-2.4642378e-008 walpha0=-1.0265377e-013 wbeta0=2.234567e-007 wint=-1e-008 wk1=6.795952e-008 wk2=-2.1981336e-008 wketa=-7.3317252e-009 wkt1=-1.1400184e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=3.0548187e-008 wtvoff=0 wu0=5.9658614e-010 wua1=1.7890568e-016 wua=-7.884629e-018 wub1=-1.3550978e-025 wub=-4.9106352e-027 wuc1=4.1267577e-017 wuc=-1.4037289e-017 wvoff=-1.6675146e-009 wvth0=4.5642665e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.1 pmos a0=1.1459651 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19108744 alpha0=7.4846555e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=42.345869 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0114756 k2=-0.018690632 k3=0 k3b=0 keta=-0.0053017786 kt1=-0.30808974 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.5959096e-007 lags=1.0404081e-007 lalpha0=-3.4131346e-011 lbeta0=-4.8401083e-006 level=54 lint=0 lk1=-6.5471375e-008 lk2=-5.6604249e-010 lketa=-2.1929041e-008 lkt1=-3.5941865e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=1.1879561e-007 lpdiblc2=2.3979675e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.1365149e-009 lua=8.3937346e-016 lub1=-5.9423465e-025 lub=-3.4811665e-025 luc1=-3.0172107e-017 luc=5.7491694e-017 lvoff=1.259976e-008 lvth0=7.848145e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.6768655e-014 pags=-3.0843241e-014 palpha0=-2.407651e-018 paramchk=1 pbeta0=8.5825341e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.25477175 pdiblc1=0.1484 pdiblc2=0.00024955823 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=2.1748834e-014 pk2=-6.129007e-015 pketa=1.1103413e-015 pkt1=-1.6287571e-014 ppclm=-2.1664163e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-9.9642066e-017 pua=-1.6983026e-022 pub1=9.6755564e-032 pub=9.5816488e-032 puc1=3.2782971e-024 puc=-7.5182999e-024 pvag=0 pvth0=1.5317707e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.01031351 ua1=1.5e-009 ua=3.8413264e-010 ub1=-2.2459185e-018 ub=1.0907567e-018 uc1=-7.622458e-011 uc=-1.2185662e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12347027 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.71729526 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=3.9893726e-008 wags=1.3857952e-008 walpha0=4.918957e-012 wbeta0=2.85852e-007 wint=-1e-008 wk1=-1.8245666e-008 wk2=-2.6841281e-009 wketa=-2.2567913e-009 wkt1=2.5589445e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=8.7678071e-008 wtvoff=0 wu0=-2.5501298e-010 wua=-4.6769074e-017 wub1=-3.2798588e-026 wub=-1.9694477e-025 wuc1=6.4565445e-018 wuc=-7.7156746e-018 wvth0=6.1706137e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.2 pmos a0=1.2624795 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.15738448 alpha0=0.0020563928 alpha1=0 at=12000 b0=0 b1=0 beta0=44.429178 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95371136 k2=-0.010397236 k3=0 k3b=0 keta=-4.2919829e-005 kt1=-0.26812521 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-3.9847608e-007 lags=1.4421474e-007 lalpha0=-2.3961345e-009 lbeta0=-7.3234127e-006 level=54 lint=0 lk1=3.3836545e-009 lk2=-1.045177e-008 lketa=-2.8197601e-008 lkt1=-5.1231914e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4138473e-007 lpclm=3.9541387e-008 lpdiblc2=4.4342116e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=3.0063094e-009 lua=8.1940101e-016 lub1=3.3763797e-025 lub=-6.8481784e-026 luc1=-7.9159583e-017 luc=9.5540362e-017 lvoff=-1.8037078e-008 lvoffcv=-2.1655389e-007 lvth0=-9.6535664e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9458182 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=3.495459e-014 pags=-1.520792e-014 palpha0=-2.3868227e-017 paramchk=1 pbeta0=-6.9013864e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32126019 pdiblc1=0.1484 pdiblc2=7.8732382e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-3.755349e-014 pk2=9.1608133e-015 pketa=2.6725774e-015 pkt1=2.6896755e-014 ppclm=7.6673781e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-6.7198364e-016 pua=-1.6075256e-022 pub1=-1.7725993e-031 pub=-4.2154414e-033 puc1=2.6039988e-023 puc=-1.8979559e-023 pvag=0 pvoff=-1.2167579e-015 pvth0=4.3646606e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0087448909 ua1=1.5e-009 ua=4.0088804e-010 ub1=-3.0276908e-018 ub=8.5616366e-019 uc1=-3.5127704e-011 uc=-4.4105686e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097768223 voffcv=0.021672727 voffl=0 vsat=94000 vth0=-0.70261262 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-3.4982576e-009 wags=7.410721e-010 walpha0=2.2922796e-011 wbeta0=4.1575066e-007 wint=-1e-008 wk1=3.1504606e-008 wk2=-1.5511159e-008 wketa=-3.567392e-009 wkt1=-1.0639016e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=5.1797956e-009 wtvoff=0 wu0=2.2513935e-010 wua=-5.4384592e-017 wub1=1.9708019e-025 wub=-1.1302537e-025 wuc1=-1.2638834e-017 wuc=1.8994754e-018 wvoff=1.0207701e-009 wvth0=3.7940282e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.3 pmos a0=1.2226 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.1718175 alpha0=0.0018165875 alpha1=0 at=12000 b0=0 b1=0 beta0=43.69625 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95405 k2=-0.01144325 k3=0 k3b=0 keta=-0.0028649375 kt1=-0.2732525 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3252175 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0090457625 ua1=1.5e-009 ua=4.8289375e-010 ub1=-2.9939e-018 ub=8.4931e-019 uc1=-4.305e-011 uc=-3.4544e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.099573375 voffcv=0 voffl=0 vsat=94000 vth0=-0.70357875 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-7.809375e-010 walpha0=2.0534062e-011 wbeta0=4.0884375e-007 wint=-1e-008 wk1=2.774625e-008 wk2=-1.4594344e-008 wketa=-3.2999203e-009 wkt1=-7.9471875e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=1.2853312e-008 wtvoff=0 wu0=1.5788719e-010 wua=-7.0472719e-017 wub1=1.7934e-025 wub=-1.1344725e-025 wuc1=-1.003275e-017 wvoff=8.9899687e-010 wvth0=4.2308437e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.4 pmos a0=0.66090759 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20881855 alpha0=1.1910101e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=38.07575 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99667836 k2=0.013187532 k3=0 k3b=0 keta=-0.10373614 kt1=-0.33233495 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-9.8161425e-008 lags=6.6568316e-008 lalpha0=-2.8926407e-012 lbeta0=-2.59284e-006 level=54 lint=0 lk1=-3.3863555e-008 lk2=-1.9573129e-008 lketa=2.1193464e-008 lkt1=5.5962764e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=2.5826511e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.7578086e-009 lua1=-2.459016e-016 lua=7.1544135e-016 lub1=-2.7023324e-026 lub=-2.9606431e-025 luc1=-3.3340425e-017 luc=1.1953068e-017 lvth0=-2.0423367e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-5.3656847e-014 pags=6.0469439e-015 palpha0=7.2099467e-020 paramchk=1 pbeta0=-3.4314451e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.37955209 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=1.0814082e-015 pketa=-3.4448579e-015 pkt1=-6.438151e-015 ppclm=2.829545e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-2.0175109e-016 pua1=1.2909834e-022 pua=-3.9456029e-023 pub1=-1.7956405e-031 pub=8.4668392e-032 puc1=3.3330844e-023 puc=-6.3347605e-024 pvag=0 pvth0=-5.0856922e-016 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0092992182 ua1=1.9998e-009 ua=-3.8099091e-011 ub1=-2.8913745e-018 ub=1.7356567e-018 uc1=5.1850909e-012 uc=8.7523896e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.70624891 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.9726782e-007 wags=-3.0445036e-008 walpha0=-4.1353238e-013 wbeta0=1.0015544e-006 wint=-1e-008 wk2=-1.3793528e-008 wketa=1.2664919e-008 wkt1=1.386661e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.9829298e-008 wtvoff=0 wu0=-1.7793682e-010 wua1=-2.62395e-016 wua=4.2158932e-017 wub1=2.6243509e-025 wub=-5.6840223e-025 wuc1=-9.3985118e-017 wuc=-1.3875714e-017 wvth0=1.5072177e-008 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.5 pmos a0=1.3400455 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19317874 alpha0=0.00012240188 alpha1=0 at=12000 b0=0 b1=0 beta0=43.297479 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.976722 k2=-0.026858767 k3=0 k3b=0 keta=-0.0020187086 kt1=-0.28407944 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-4.3229728e-007 lags=7.4263098e-008 lalpha0=-5.7254595e-011 lbeta0=-5.1619305e-006 level=54 lint=0 lk1=-2.4045024e-008 lk2=1.2965043e-010 lketa=-2.8851515e-008 lkt1=-2.3182084e-008 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=-5.9115571e-008 lpdiblc2=2.3979675e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.5273198e-009 lua=5.6122091e-016 lub1=9.5153784e-026 lub=-6.9209035e-026 luc1=1.7945798e-017 luc=5.0666426e-017 lvoff=1.259976e-008 lvth0=-3.6235097e-010 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.3902161e-014 pags=-1.5209944e-014 palpha0=9.7320549e-018 paramchk=1 pbeta0=2.5478195e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.5521986 pdiblc1=0.1484 pdiblc2=0.00024955823 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-6.4942458e-015 pketa=4.7446404e-015 pkt1=-6.0039252e-015 ppclm=7.1739209e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-3.0481466e-016 pua=-2.3800175e-023 pub1=-2.6517336e-031 pub=-5.0610011e-032 puc1=-2.1983603e-023 puc=-3.9350342e-024 pvag=0 pvth0=5.8422811e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097676914 ua1=1.5e-009 ua=2.7535709e-010 ub1=-3.139702e-018 ub=1.2745688e-018 uc1=-9.90552e-011 uc=8.8382089e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12347027 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.70966351 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-6.1998457e-008 wags=1.276002e-008 walpha0=-2.0047588e-011 wbeta0=-2.1374325e-007 wint=-1e-008 wk2=1.6041428e-009 wketa=-3.980403e-009 wkt1=1.2984037e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-6.8471025e-008 wtvoff=0 wu0=3.1542e-011 wua=1.033809e-017 wub1=4.3643775e-025 wub=-2.9344612e-025 wuc1=1.844262e-017 wuc=-1.8753207e-017 wvth0=2.163945e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.6 pmos a0=1.1183126 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16571096 alpha0=0.0021722983 alpha1=0 at=12000 b0=0 b1=0 beta0=44.346784 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0137201 k2=-0.027400332 k3=0 k3b=0 keta=-0.0068379523 kt1=-0.33792326 kt1l=0 kt2=-0.016960609 ku0=0 kvsat=0 kvth0=0 la0=-1.6799168e-007 lags=1.0700469e-007 lalpha0=-2.5007312e-009 lbeta0=-6.4127021e-006 level=54 lint=0 lk1=-6.8146803e-008 lk2=7.7519526e-010 lketa=-2.3106977e-008 lkt1=4.0999742e-008 lkt2=4.642374e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4138473e-007 lpclm=2.0695108e-007 lpdiblc2=4.4342116e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.5655154e-009 lua=4.0804167e-016 lub1=-5.516372e-025 lub=5.7383397e-026 luc1=-4.9455495e-017 luc=5.9563621e-017 lvoff=-2.0354712e-008 lvoffcv=-2.1655389e-007 lvth0=-1.3636128e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9458182 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-8.6049719e-014 pags=4.3273558e-015 palpha0=3.1045047e-017 paramchk=1 pbeta0=-5.4713694e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32898832 pdiblc1=0.1484 pdiblc2=7.8732382e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=3.2666562e-015 pkt1=-2.1524865e-014 pkt2=-2.4372464e-015 ppclm=-1.1216307e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=8.4433178e-017 pua=5.5211091e-023 pub1=2.8960953e-031 pub=-7.0294662e-032 puc1=1.0445342e-023 puc=-9.1769787e-026 pvag=0 pvth0=1.2434931e-017 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097356481 ua1=1.5e-009 ua=4.0386316e-010 ub1=-2.5970921e-018 ub=1.1683671e-018 uc1=-4.2510491e-011 uc=1.3741189e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.095823899 voffcv=0.021672727 voffl=0 vsat=94000 vth0=-0.70882353 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=7.2189361e-008 wags=-3.630332e-009 walpha0=-3.7927615e-011 wbeta0=4.590075e-007 wint=-1e-008 wk2=-6.5845334e-009 wkt1=2.600496e-008 wkt2=2.0446698e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.1225287e-009 wtvoff=0 wu0=-2.950082e-010 wua=-5.594653e-017 wub1=-2.898414e-026 wub=-2.7693216e-025 wuc1=-8.7628704e-018 wuc=-2.1977422e-017 wvth0=7.0547555e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.7 pmos a0=1.1015 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17642 alpha0=0.001922025 alpha1=0 at=12000 b0=0 b1=0 beta0=43.705 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.02732275 k3=0 k3b=0 keta=-0.0091505 kt1=-0.33382 kt1l=0 kt2=-0.016496 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.009892325 ua1=1.5e-009 ua=4.447e-010 ub1=-2.6523e-018 ub=1.17411e-018 uc1=-4.746e-011 uc=7.33525e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0=-0.70896 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=6.35775e-008 wags=-3.19725e-009 walpha0=-3.4820625e-011 wbeta0=4.0425e-007 wint=-1e-008 wk2=-6.2576062e-009 wkt1=2.385075e-008 wkt2=1.80075e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wtvoff=0 wu0=-2.8655813e-010 wua=-5.0421e-017 wub=-2.8396725e-025 wuc1=-7.7175e-018 wuc=-2.1986606e-017 wvth0=7.056e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.8 pmos a0=0.87958485 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.33412256 alpha0=9.5916748e-006 alpha1=0 at=12000 b0=0 b1=0 beta0=37.669715 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99667836 k2=-0.0016908531 k3=0 k3b=0 keta=-0.087907195 kt1=-0.29643476 kt1l=0 kt2=-0.020721765 ku0=0 kvsat=0 kvth0=0 la0=-1.4075717e-007 lags=-2.3726975e-009 lalpha0=-2.1820478e-012 lbeta0=-2.2686901e-006 level=54 lint=0 lk1=-3.3863555e-008 lk2=-1.6910112e-008 lketa=1.6887989e-008 lkt1=-8.0291808e-009 lkt2=2.0823681e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=4.8328885e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.7102254e-009 lua1=-1.4896941e-016 lua=6.0284809e-016 lub1=-1.2288098e-025 lub=3.159209e-026 luc1=8.5354274e-019 luc=-7.1184051e-018 lvth0=-8.3892994e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.4770608e-015 pags=9.0499685e-014 palpha0=-7.9837683e-019 paramchk=1 pbeta0=-7.4022817e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32767553 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-2.1807869e-015 pketa=1.8293483e-015 pkt1=4.0831393e-015 pkt2=-2.550901e-015 ppclm=7.3004154e-016 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.4346165e-016 pua1=1.0356403e-023 pua=9.847072e-023 pub1=-6.213842e-032 pub=-3.167107e-031 puc1=-8.556766e-024 puc=1.7027795e-023 pvag=0 pvth0=7.26646e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011456358 ua1=1.8027834e-009 ua=3.841223e-010 ub1=-2.5917035e-018 ub=9.2943227e-019 uc1=-8.5734843e-011 uc=1.3336117e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.69776909 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-7.0611818e-008 wags=-1.8394245e-007 walpha0=2.4265399e-012 wbeta0=1.4989467e-006 wint=-1e-008 wk2=4.4324937e-009 wketa=-6.7255452e-009 wkt1=-3.0111128e-008 wkt2=9.3783124e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=8.3378086e-008 wtvoff=0 wu0=-2.8204333e-009 wua1=-2.10496e-017 wua=-4.7506228e-016 wub1=-1.0466188e-025 wub=4.1922273e-025 wuc1=1.7391801e-017 wuc=-7.0026382e-017 wvth0=4.6843987e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.9 pmos a0=1.1742768 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20869703 alpha0=0.00011037751 alpha1=0 at=12000 b0=0 b1=0 beta0=43.119792 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.976722 k2=-0.03059107 k3=0 k3b=0 keta=-0.0069935214 kt1=-0.3027753 kt1l=0 kt2=-0.010659902 ku0=0 kvsat=0 kvth0=0 la0=-2.8574559e-007 lags=5.9336662e-008 lalpha0=-5.1768678e-011 lbeta0=-4.9501275e-006 level=54 lint=0 lk1=-2.4045024e-008 lk2=-2.6912057e-009 lketa=-2.2921538e-008 lkt1=-4.9096367e-009 lkt2=-2.8680684e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.3546458e-008 lpdiblc2=2.3979675e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.3484099e-009 lua=6.2730931e-016 lub1=-1.8564299e-025 lub=1.538535e-026 luc1=-2.4051688e-017 luc=7.1676685e-017 lvoff=-1.7539439e-009 lvth0=-6.989061e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.0562366e-013 pags=3.0749415e-015 palpha0=3.0118059e-018 paramchk=1 pbeta0=-4.6767172e-015 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.37804632 pdiblc1=0.1484 pdiblc2=0.00024955823 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-3.038697e-015 pketa=-2.5195814e-015 pkt1=-2.8387673e-014 pkt2=3.5133838e-015 ppclm=-2.9521777e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.31065e-015 pua=-1.0475847e-022 pub1=7.8802685e-032 pub=-1.5423813e-031 puc1=2.9463318e-023 puc=-2.9672601e-023 pvag=0 pvoff=1.7583287e-014 pvth0=1.3960001e-014 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010159235 ua1=1.5e-009 ua=3.3440437e-010 ub1=-2.4641385e-018 ub=9.623728e-019 uc1=-3.5114455e-011 uc=-2.6791447e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094296073 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.7006151 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.4106826e-007 wags=-6.2498812e-009 walpha0=-5.3177339e-012 wbeta0=3.9234204e-009 wint=-1e-008 wk2=6.1762134e-009 wketa=2.1137428e-009 wkt1=3.5886458e-008 wkt2=-2.9474696e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.4486552e-007 wtvoff=0 wu0=-4.4809927e-010 wua=-6.1994828e-017 wub1=-3.9112754e-025 wub=8.8993941e-026 wuc1=-5.9884793e-017 wuc=2.4893122e-017 wvoff=-3.5738389e-008 wvth0=-8.9203589e-009 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.10 pmos a0=1.1830432 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16693357 alpha0=0.0021410284 alpha1=0 at=12000 b0=0 b1=0 beta0=44.157511 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0137201 k2=-0.03602212 k3=0 k3b=0 keta=-0.0068379523 kt1=-0.29670745 kt1l=0 kt2=-0.012756202 ku0=0 kvsat=0 kvth0=0 la0=-2.9619524e-007 lags=1.0911871e-007 lalpha0=-2.4723045e-009 lbeta0=-6.1870892e-006 level=54 lint=0 lk1=-6.8146803e-008 lk2=3.7826066e-009 lketa=-2.3106977e-008 lkt1=-1.2142514e-008 lkt2=-3.6927975e-010 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4138473e-007 lpclm=6.510159e-008 lpdiblc2=4.4342116e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.306639e-009 lua1=1.2396634e-016 lua=2.2975668e-016 lub1=4.3880232e-026 luc1=1.3468483e-017 luc=5.9488707e-017 lvoff=2.8334685e-009 lvoffcv=-2.1655389e-007 lvth0=-4.4372015e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9458182 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.0999638e-014 pags=1.7376873e-015 palpha0=-3.7775811e-018 paramchk=1 pbeta0=-8.2351269e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34318463 pdiblc1=0.1484 pdiblc2=7.8732382e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-4.1742272e-016 pkt1=4.3574398e-014 pkt2=3.7020295e-015 ppclm=1.6254932e-013 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=4.0155688e-016 pua1=-1.5185876e-022 pua=2.736102e-022 pub1=-4.3989932e-031 puc1=-6.6636531e-023 pvag=0 pvoff=-2.8405521e-014 pvth0=3.7775811e-015 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011033204 ua1=1.3960014e-009 ua=6.6792168e-010 ub1=-2.6566915e-018 ub=9.7527997e-019 uc1=-6.6591108e-011 uc=-1.6566634e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.098144574 voffcv=0.021672727 voffl=0 vsat=94000 vth0=-0.70275593 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-7.1056483e-009 wags=-5.1280236e-009 walpha0=3.7806056e-013 wbeta0=6.9086635e-007 wint=-1e-008 wk2=3.9771578e-009 wkt1=-2.4484407e-008 wkt2=-3.1057295e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=-1.6267946e-008 wtvoff=0 wu0=-1.8845144e-009 wua1=1.2739829e-016 wua=-3.7941821e-016 wub1=4.4025153e-026 wub=-4.0400465e-026 wuc1=2.0735886e-017 wvoff=2.8428264e-009 wvth0=-3.7806056e-010 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.11 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17785418 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.538307 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035643557 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29792267 kt1l=0 kt2=-0.012793159 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011163973 ua1=1.4084079e-009 ua=6.9091574e-010 ub1=-2.6523e-018 ub=9.7527997e-019 uc1=-6.5243182e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0=-0.7032 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-4.9541158e-009 wbeta0=6.0844915e-007 wint=-1e-008 wk2=3.9353821e-009 wkt1=-2.0123479e-008 wkt2=-2.7352301e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wtvoff=0 wu0=-1.8443266e-009 wua1=1.1220026e-016 wua=-3.5203528e-016 wub=-4.0400465e-026 wuc1=1.4066898e-017 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.12 pmos a0=0.87254127 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.31577418 alpha0=9.8337236e-006 alpha1=0 at=12000 b0=0 b1=0 beta0=37.819236 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99667836 k2=-0.0012487091 k3=0 k3b=0 keta=-0.088578073 kt1=-0.29943836 kt1l=0 kt2=-0.019786273 ku0=0 kvsat=0 kvth0=0 la0=-1.4090451e-007 lags=6.6547025e-009 lalpha0=-2.2616864e-012 lbeta0=-2.3425283e-006 level=54 lint=0 lk1=-3.3863555e-008 lk2=-1.7127647e-008 lketa=1.7070468e-008 lkt1=-7.6218851e-009 lkt2=1.8279142e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=4.8401708e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.695915e-009 lua1=-1.4793635e-016 lua=6.126706e-016 lub1=-1.2907933e-025 luc=-5.419872e-018 lvth0=-7.6644654e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.33599254 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011175018 ua1=1.8006836e-009 ua=3.3673455e-010 ub1=-2.6021436e-018 ub=9.7125e-019 uc1=-8.4e-011 uc=1.26376e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.69730182 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.13 pmos a0=1.1883484 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.2080736 alpha0=0.00010984706 alpha1=0 at=12000 b0=0 b1=0 beta0=43.120183 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.976722 k2=-0.029974989 k3=0 k3b=0 keta=-0.0067826743 kt1=-0.2991956 kt1l=0 kt2=-0.010953914 ku0=0 kvsat=0 kvth0=0 la0=-2.9628161e-007 lags=5.9643389e-008 lalpha0=-5.1468248e-011 lbeta0=-4.950594e-006 level=54 lint=0 lk1=-2.4045024e-008 lk2=-2.9943176e-009 lketa=-2.3172868e-008 lkt1=-7.7413248e-009 lkt2=-2.5176062e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.0601642e-008 lpdiblc2=2.3979675e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.2176717e-009 lua=6.1685959e-016 lub1=-1.7778237e-025 luc1=-2.1112704e-017 luc=6.8716825e-017 lvth0=-5.5965422e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.39249674 pdiblc1=0.1484 pdiblc2=0.00024955823 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010114537 ua1=1.5e-009 ua=3.2822034e-010 ub1=-2.5031537e-018 ub=9.7125e-019 uc1=-4.1088e-011 uc=-2.4308343e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0=-0.70150491 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.14 pmos a0=1.1823344 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16642204 alpha0=0.0021410661 alpha1=0 at=12000 b0=0 b1=0 beta0=44.226425 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0137201 k2=-0.035625396 k3=0 k3b=0 keta=-0.0068379523 kt1=-0.29914978 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.8911298e-007 lags=1.0929204e-007 lalpha0=-2.4726813e-009 lbeta0=-6.2692351e-006 level=54 lint=0 lk1=-6.8146803e-008 lk2=3.7409685e-009 lketa=-2.3106977e-008 lkt1=-7.7959401e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4138473e-007 lpclm=8.1315986e-008 lpdiblc2=4.4342116e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.3466945e-009 lua1=1.0881833e-016 lua=2.5704947e-016 luc1=6.8214476e-018 luc=5.9488707e-017 lvoffcv=-2.1655389e-007 lvth0=-4.0603855e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9458182 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34156189 pdiblc1=0.1484 pdiblc2=7.8732382e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010845223 ua1=1.4087095e-009 ua=6.3007447e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.4522691e-011 uc=-1.6566634e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0.021672727 voffl=0 vsat=94000 vth0=-0.70279364 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.model pmos_3p3.15 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17736 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.599 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=3.8e-011 cgdo=1.178e-010 cgidl=7.5 cgsl=3.8e-011 cgso=1.178e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035251 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29993 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw=466 rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe=7.7e-009 toxm=7.9e-009 toxp=7.7e-009 toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.01098 ua1=1.4196e-009 ua=6.558e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.384e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0=-0.7032 vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj=1e-007 xl=-8e-009 xpart=0 xtis=3 xw=5e-009
.subckt pplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 par=1 r_rsh0='rsh_pplus_u_m' r_dw=2.75e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.375e-3 r_tc2=1e-6 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model pn_junction d cj=0.00094344 level=2
d1 1 3 pn_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends pplus_u_m1
.endl pmos_3p3_sf

.lib nmos_6p0_t
.subckt nmos_6p0_sab d g s b w=10u l=0.6u par=1 s_sab=0.28u d_sab=3.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.01155
.param par_k=0.0000
.param par_l=4e-7
.param par_w=-5e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b nplus_u_m2 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b nplus_u_m2 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b nmos_6p0 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='0' sb='0' sd='0' delvto='mis_vth*sw_stat_mismatch'
.ends
.model nmos_6p0.0 nmos a0=0.72499969 a1=0 a2=0.96 acde=0.3 acnqsmod=0 agidl=0 ags=0.13699995 aigbacc=0.43 aigbinv=0.35 aigc=0.43 aigsd=0.43 alpha0=-1.88e-007 alpha1=19 at=109000.03 b0=0 b1=0 beta0=36.6 bgidl=2.3e+009 bigbacc=0.054 bigbinv=0.03 bigc=0.054 bigsd=0.054 binunit=1 bvs=11 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cgbo=1e-013 cgdl='1.5e-010*nmos_6p0_cgdo' cgdo='1e-010*nmos_6p0_cgdo' cgidl=0.5 cgsl='1.5e-010*nmos_6p0_cgso' cgso='1e-010*nmos_6p0_cgso' cigbacc=0.075 cigbinv=0.006 cigc=0.075 cigsd=0.075 cit=0 cjs=0.00095 cjswgs=3.573e-010 cjsws=1.33e-010 ckappad=0.6 ckappas=0.6 clc=1e-010 cle=0.6 delta=0.01 diomod=1 dlc=5.4e-8 dlcig=0 dmcg=0 dmcgt=0 dmdg=0 drout=0.4 dsub=0.4 dvt0=5.72 dvt0w=10 dvt1=0.299 dvt1w=976700 dvt2=-0.0793 dvt2w=0.15 dvtp0=0 dvtp1=0 dwb=6e-009 dwc=0 dwg=-6e-010 ef=1 egidl=0.8 eigbinv=1.1 em=4.1e+007 epsrox=3.9 eta0=0 etab=-0.43 eu=1.67 fnoimod=1 fprout=0 gbmin=1e-012 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=6.88e-007 jswgs=0 jsws=4.88e-013 jtsd=0 jtss=0 jtsswd=0 jtsswgd=0 jtsswgs=0 jtssws=0 k1=0.9 k2=-0.001 k2we=0 k3=-1.1369995 k3b=0.86 keta=-0.021200021 kt1=-0.412 kt1l=3.5e-008 kt2=-0.05 ku0=0 ku0we=0 kvsat=0 kvth0=0 kvth0we=0 la0=0.40144032 lags=-0.068999933 lambda=0 lat=-75600.021 level=54 lint=-3e-008 lintnoi=0 lketa=0.04140001 lku0=0 lkvth0=0 ll=1.93e-014 llc=0 lln=1 llodku0=0 llodvth=0 lmax=5.0001e-005 lmin=7e-007 lodeta0=1 lodk2=1 lp=1e-008 lpclm=0.89088024 lpe0=1.63e-007 lpeb=0 lu0=0.019999998 lua=-3.3696895e-019 lub=1.7400001e-018 luc1=-1.8816003e-011 luc=9.8000018e-011 lute=0.030000222 lvsat='-2649.9871*nmos_6p0_vsat' lw=0 lwc=0 lwl=0 lwlc=0 lwn=1 minv=0 mjs=0.296 mjswgs=0.40313 mjsws=0.01 mobmod=0 moin=15 ndep=1.7e+017 nfactor=0.864 ngate=1e+020 ngcon=1 nigbacc=1 nigbinv=3 nigc=1 njs=1.0541 njts=20 njtssw=20 njtsswg=20 noff=1.5 noia='nmos_6p0_noia' noib='nmos_6p0_noib' noic='nmos_6p0_noic' nsd=1e+020 ntnoi=1 ntox=1 pags=0.0070910278 paramchk=1 pat=-6699.9857 pbs=0.606 pbswgs=0.861 pbsws=0.48 pclm=0.0099999763 pdiblc1=1.6 pdiblc2=0.0022 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pigcd=1 pku0=0 pkvth0=0 poxedge=1 prt=0 prwb=0 prwg=1 pscbe1=4.325e+009 pscbe2=8.8e-006 pu0=0.0018000065 pua=1.4622721e-010 pub=-2.3803999e-019 puc=-5.6168065e-012 pute=-0.019999981 pvag=1.75 pvsat='6308.7992*nmos_6p0_vsat' rbdb=50 rbdbx0=100 rbdby0=100 rbodymod=0 rbpb=50 rbpbx0=100 rbpbxl=0 rbpbxnf=0 rbpbxw=0 rbpby0=100 rbpbyl=0 rbpbynf=0 rbpbyw=0 rbpd0=50 rbpd=50 rbpdl=0 rbpdnf=0 rbpdw=0 rbps0=50 rbps=50 rbpsl=0 rbpsnf=0 rbpsw=0 rbsb=50 rbsbx0=100 rbsby0=100 rbsdbxl=0 rbsdbxnf=0 rbsdbxw=0 rbsdbyl=0 rbsdbynf=0 rbsdbyw=0 rdsmod=0 rdsw=2175 rdswmin=0 rdw=100 rdwmin=0 rgatemod=0 rsh=7 rshg=0.1 rsw=100 rswmin=0 saref=1e-006 sbref=1e-006 scref=1e-006 steta0=0 stk2=0 tcj=0.000825 tcjsw=0.0018 tcjswg=0.001595 tempmod=0 tku0=0 tnjts=0 tnjtssw=0 tnjtsswg=0 tnoimod=0 tnom=25 toxe='1.52e-008+nmos_6p0_tox' toxm='1.52e-008+nmos_6p0_tox' toxp='1.6e-008+nmos_6p0_tox' toxref=1.52e-008 tpb=0.00146 tpbsw=0.00313 tpbswg=0.0016588 trnqsmod=0 tvfbsdoff=0 tvoff=0 u0=0.052500014 ua1=1e-009 ua=6.8000001e-012 ub1=-1e-018 ub=2.8799997e-018 uc1=-5.5999995e-011 uc=7.9399996e-011 ud1=0 up=0 ute=-1.5000005 vbm=-3 version=4.5 vfbcv=-1 vfbsdoff=0 voff=-0.08 voffcv=0 voffl=0 vsat='103999.98*nmos_6p0_vsat' vth0='0.67314+nmos_6p0_vth0' vtl=200000 vtsd=10 vtss=10 vtsswd=10 vtsswgd=10 vtsswgs=10 vtssws=10 w0=1e-009 wags=-4.2211594e-008 wat=6479.9797 web=0 wec=0 wint=1.55e-008 wk3=-0.047531062 wku0=0 wkvth0=0 wl=0 wlc=0 wln=1 wlod=0 wlodku0=0 wlodvth=0 wmax=0.000100001 wmin=3e-007 wpemod=0 wr=1 wu0=-8.0300635e-009 wua=-8.4912706e-019 wub=-1.1655759e-026 wuc=8.0000028e-012 wute=0.06000001 wvsat='0.012447116*nmos_6p0_vsat' ww=-2.7e-015 wwc=0 wwl=0 wwlc=0 wwn=1 xgl=0 xgw=0 xj=1.5e-007 xjbvd=1 xjbvs=1 xl='0+nmos_6p0_xl' xn=3 xpart=0 xrcrg1=12 xrcrg2=1 xtis=3 xtsd=0.02 xtss=0.02 xtsswd=0.02 xtsswgd=0.02 xtsswgs=0.02 xtssws=0.02 xw='0+nmos_6p0_xw'
.model nmos_6p0.1 nmos a0=0.72500081 a1=0 a2=0.96 acde=0.3 acnqsmod=0 agidl=0 ags=0.13700019 aigbacc=0.43 aigbinv=0.35 aigc=0.43 aigsd=0.43 alpha0=-1.88e-007 alpha1=19 at=-119957.68 b0=0 b1=0 beta0=36.6 bgidl=2.3e+009 bigbacc=0.054 bigbinv=0.03 bigc=0.054 bigsd=0.054 binunit=1 bvs=11 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cgbo=1e-013 cgdl='1.5e-010*nmos_6p0_cgdo' cgdo='1e-010*nmos_6p0_cgdo' cgidl=0.5 cgsl='1.5e-010*nmos_6p0_cgso' cgso='1e-010*nmos_6p0_cgso' cigbacc=0.075 cigbinv=0.006 cigc=0.075 cigsd=0.075 cit=0 cjs=0.00095 cjswgs=3.573e-010 cjsws=1.33e-010 ckappad=0.6 ckappas=0.6 clc=1e-010 cle=0.6 delta=0.01 diomod=1 dlc=5.4e-8 dlcig=0 dmcg=0 dmcgt=0 dmdg=0 drout=0.4 dsub=0.4 dvt0=5.72 dvt0w=10 dvt1=0.299 dvt1w=976700 dvt2=-0.0793 dvt2w=0.15 dvtp0=0 dvtp1=0 dwb=6e-009 dwc=0 dwg=-6e-010 ef=1 egidl=0.8 eigbinv=1.1 em=4.1e+007 epsrox=3.9 eta0=0 etab=-0.43 eu=1.67 fnoimod=1 fprout=0 gbmin=1e-012 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=6.88e-007 jswgs=0 jsws=4.88e-013 jtsd=0 jtss=0 jtsswd=0 jtsswgd=0 jtsswgs=0 jtssws=0 k1=0.9 k2=-0.001 k2we=0 k3=-1.1369995 k3b=0.86 keta=-0.021200265 kt1=-0.412 kt1l=3.5e-008 kt2=-0.05 ku0=0 ku0we=0 kvsat=0 kvth0=0 kvth0we=0 la0=0.40143954 lags=-0.069000099 lambda=0 lat=85782.454 level=54 lint=-3e-008 lintnoi=0 lketa=0.041400183 lku0=0 lkvth0=0 ll=1.93e-014 llc=0 lln=1 llodku0=0 llodvth=0 lmax=7e-007 lmin=6e-007 lodeta0=1 lodk2=1 lp=1e-008 lpclm=0.89088046 lpe0=1.63e-007 lpeb=0 lu0=0.019999754 lua=3.7339196e-019 lub=1.7399991e-018 luc1=-1.8816017e-011 luc=9.7999741e-011 lute=0.030000412 lvsat='24946.5*nmos_6p0_vsat' lw=0 lwc=0 lwl=0 lwlc=0 lwn=1 minv=0 mjs=0.296 mjswgs=0.40313 mjsws=0.01 mobmod=0 moin=15 ndep=1.7e+017 nfactor=0.864 ngate=1e+020 ngcon=1 nigbacc=1 nigbinv=3 nigc=1 njs=1.0541 njts=20 njtssw=20 njtsswg=20 noff=1.5 noia='nmos_6p0_noia' noib='nmos_6p0_noib' noic='nmos_6p0_noic' nsd=1e+020 ntnoi=1 ntox=1 pags=0.0070909573 paramchk=1 pat=21832.424 pbs=0.606 pbswgs=0.861 pbsws=0.48 pclm=0.0099996572 pdiblc1=1.6 pdiblc2=0.0022 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pigcd=1 pku0=0 pkvth0=0 poxedge=1 prt=0 prwb=0 prwg=1 pscbe1=4.325e+009 pscbe2=8.8e-006 pu0=0.0018000207 pua=1.4622711e-010 pub=-2.3804013e-019 puc=-5.6167642e-012 pute=-0.020000108 pvag=1.75 pvsat='6308.7053*nmos_6p0_vsat' rbdb=50 rbdbx0=100 rbdby0=100 rbodymod=0 rbpb=50 rbpbx0=100 rbpbxl=0 rbpbxnf=0 rbpbxw=0 rbpby0=100 rbpbyl=0 rbpbynf=0 rbpbyw=0 rbpd0=50 rbpd=50 rbpdl=0 rbpdnf=0 rbpdw=0 rbps0=50 rbps=50 rbpsl=0 rbpsnf=0 rbpsw=0 rbsb=50 rbsbx0=100 rbsby0=100 rbsdbxl=0 rbsdbxnf=0 rbsdbxw=0 rbsdbyl=0 rbsdbynf=0 rbsdbyw=0 rdsmod=0 rdsw=2175 rdswmin=0 rdw=100 rdwmin=0 rgatemod=0 rsh=7 rshg=0.1 rsw=100 rswmin=0 saref=1e-006 sbref=1e-006 scref=1e-006 steta0=0 stk2=0 tcj=0.000825 tcjsw=0.0018 tcjswg=0.001595 tempmod=0 tku0=0 tnjts=0 tnjtssw=0 tnjtsswg=0 tnoimod=0 tnom=25 toxe='1.52e-008+nmos_6p0_tox' toxm='1.52e-008+nmos_6p0_tox' toxp='1.6e-008+nmos_6p0_tox' toxref=1.52e-008 tpb=0.00146 tpbsw=0.00313 tpbswg=0.0016588 trnqsmod=0 tvfbsdoff=0 tvoff=0 u0=0.052500361 ua1=1e-009 ua=6.7999991e-012 ub1=-1e-018 ub=2.8800011e-018 uc1=-5.5999975e-011 uc=7.9400388e-011 ud1=0 up=0 ute=-1.5000008 vbm=-3 version=4.5 vfbcv=-1 vfbsdoff=0 voff=-0.08 voffcv=0 voffl=0 vsat='64848.09*nmos_6p0_vsat' vth0='0.67314+nmos_6p0_vth0' vtl=200000 vtsd=10 vtss=10 vtsswd=10 vtsswgd=10 vtsswgs=10 vtssws=10 w0=1e-009 wags=5.7853969e-008 wat=-33999.727 web=0 wec=0 wint=1.55e-008 wk3=-0.047531062 wku0=0 wkvth0=0 wl=0 wlc=0 wln=1 wlod=0 wlodku0=0 wlodvth=0 wmax=0.000100001 wmin=3e-007 wpemod=0 wr=1 wu0=-2.8167565e-008 wua=1.3244868e-016 wub=1.8765824e-025 wuc=7.9999428e-012 wute=0.060000189 wvsat='0.14568305*nmos_6p0_vsat' ww=-2.7e-015 wwc=0 wwl=0 wwlc=0 wwn=1 xgl=0 xgw=0 xj=1.5e-007 xjbvd=1 xjbvs=1 xl='0+nmos_6p0_xl' xn=3 xpart=0 xrcrg1=12 xrcrg2=1 xtis=3 xtsd=0.02 xtss=0.02 xtsswd=0.02 xtsswgd=0.02 xtsswgs=0.02 xtssws=0.02 xw='0+nmos_6p0_xw'
.subckt nplus_u_m2 1 2 3 r_length='lr' r_width='wr' dtemp=0 r_rsh0='rsh_nplus_u_m' r_dw=-5e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.36e-3 r_tc2=6.5e-7 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model np_junction d cj=0.00096797 level=2
d1 3 1 np_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends nplus_u_m2
.endl nmos_6p0_t

.lib nmos_6p0_nat_t
.subckt nmos_6p0_nat d g s b w=1e-5 l=1.8e-6 as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 par=1 dtemp=0 sa=0 sb=0 nf=1 sd=0 m=1
m0 d g s b nmos_6p0_nat m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' sa='sa' sb='sb' nf='nf' sd='sd'
.ends nmos_6p0_nat
.model nmos_6p0_nat.0 nmos a0=0.88 a1=0 a2=0.47 acde=0.3 acnqsmod=0 agidl=2e-010 ags=0.72 aigbacc=0.43 aigbinv=0.35 aigc=0.43 aigsd=0.43 alpha0=1.36e-008 alpha1=1e-005 at=80000 b0=3.5e-007 b1=0 beta0=15 bgidl=2.3e+009 bigbacc=0.054 bigbinv=0.03 bigc=0.054 bigsd=0.054 binunit=1 bvs=11 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cgbo=1e-013 cgdl=1.5e-010 cgdo='nmos_6p0_nat_cgdo' cgidl=0.5 cgsl=1.5e-010 cgso='nmos_6p0_nat_cgso' cigbacc=0.075 cigbinv=0.006 cigc=0.075 cigsd=0.075 cit=0 cjs=0.00095 cjswgs=3.573e-010 cjsws=1.33e-010 ckappad=0.6 ckappas=0.6 clc=1e-010 cle=0.6 delta=0.005 diomod=1 dlc=0 dlcig=0 dmcg=0 dmcgt=0 dmdg=0 drout=0.16 dsub=0.4 dvt0=2.2 dvt0w=0 dvt1=0.53 dvt1w=5300000 dvt2=-0.032 dvt2w=-0.032 dvtp0=1e-008 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1 egidl=0.8 eigbinv=1.1 em=4.1e+007 epsrox=3.9 eta0=0.06 etab=-0.43 eu=1.67 fnoimod=1 fprout=65 gbmin=1e-012 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=6.88e-007 jswgs=0 jsws=4.88e-013 jtsd=0 jtss=0 jtsswd=0 jtsswgd=0 jtsswgs=0 jtssws=0 k1=0.165 k2=-0.001 k2we=0 k3=-0.6 k3b=-0.6 keta=-0.04 kt1=-0.412 kt1l=3.5e-008 kt2=-0.05 ku0=0 ku0we=0 kvsat=0 kvth0=0 kvth0we=0 lambda=0 lat=-30000 level=54 lint=1e-007 lintnoi=0 lku0=0 lkvth0=0 ll=0 llc=0 lln=1 llodku0=0 llodvth=0 lmax=50.01e-6 lmin=1.8e-6 lnfactor=0.45 lodeta0=1 lodk2=1 lp=1e-008 lpe0=1e-007 lpeb=0 lu0=0.042 lub=3.65e-018 lute=-0.26 lvth0=-0.088 lw=0 lwc=0 lwl=0 lwlc=0 lwn=1 minv=-0.5 mjs=0.296 mjswgs=0.40313 mjsws=0.01 mobmod=0 moin=15 ndep=1.7e+017 nfactor=0.40241 ngate=1e+020 ngcon=1 nigbacc=1 nigbinv=3 nigc=1 njs=1.0541 njts=20 njtssw=20 njtsswg=20 noff=1.5 noia='nmos_6p0_nat_noia' noib='nmos_6p0_nat_noib' noic='nmos_6p0_nat_noic' nsd=1e+020 ntnoi=1 ntox=1 paramchk=1 pat=-10000 pbs=0.606 pbswgs=0.861 pbsws=0.48 pclm=3 pdiblc1=1.41 pdiblc2=1e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.5 pigcd=1 pku0=0 pkvth0=0 poxedge=1 prt=0 prwb=0 prwg=1 pscbe1=5e+009 pscbe2=5e-006 pvag=1 pvsat=23500 rbdb=50 rbdbx0=100 rbdby0=100 rbodymod=0 rbpb=50 rbpbx0=100 rbpbxl=0 rbpbxnf=0 rbpbxw=0 rbpby0=100 rbpbyl=0 rbpbynf=0 rbpbyw=0 rbpd0=50 rbpd=50 rbpdl=0 rbpdnf=0 rbpdw=0 rbps0=50 rbps=50 rbpsl=0 rbpsnf=0 rbpsw=0 rbsb=50 rbsbx0=100 rbsby0=100 rbsdbxl=0 rbsdbxnf=0 rbsdbxw=0 rbsdbyl=0 rbsdbynf=0 rbsdbyw=0 rdsmod=0 rdsw=3480 rdswmin=0 rdw=100 rdwmin=0 rgatemod=0 rsh=7 rshg=0.1 rsw=100 rswmin=0 saref=1e-006 sbref=1e-006 scref=1e-006 steta0=0 stk2=0 tcj=0.000825 tcjsw=0.0018 tcjswg=0.001595 tempmod=0 tku0=0 tnjts=0 tnjtssw=0 tnjtsswg=0 tnoimod=0 tnom=25 toxe='nmos_6p0_nat_tox' toxm=1.52e-008 toxp=1.6e-008 toxref=1.52e-008 tpb=0.00146 tpbsw=0.00313 tpbswg=0.0016588 trnqsmod=0 tvfbsdoff=0 tvoff=0 u0='nmos_6p0_nat_u0' ua1=1e-009 ua=2.278e-009 ub1=-1e-018 ub=3.97e-019 uc1=-5.6e-011 uc=2.625e-012 ud1=0 up=0 ute=-1.5 vbm=-3 version=4.5 vfbcv=-1 vfbsdoff=0 voff=-0.06 voffcv=0 voffl=0 vsat=106700 vth0='nmos_6p0_nat_vth0' vtl=200000 vtsd=10 vtss=10 vtsswd=10 vtsswgd=10 vtsswgs=10 vtssws=10 w0=1e-010 web=0 wec=0 wint=1e-009 wku0=0 wkvth0=0 wl=0 wlc=0 wln=1 wlod=0 wlodku0=0 wlodvth=0 wmax=100.01e-6 wmin=0.8e-6 wpemod=0 wr=1 ww=0 wwc=0 wwl=0 wwlc=0 wwn=1 xgl=0 xgw=0 xj=1.5e-007 xjbvd=1 xjbvs=1 xl='nmos_6p0_nat_xl' xn=3 xpart=0 xrcrg1=12 xrcrg2=1 xtis=3 xtsd=0.02 xtss=0.02 xtsswd=0.02 xtsswgd=0.02 xtsswgs=0.02 xtssws=0.02 xw='nmos_6p0_nat_xw'
.endl nmos_6p0_nat_t

.lib pmos_6p0_t
.subckt pmos_6p0_sab d g s b w=10u l=0.5u par=1 s_sab=0.28u d_sab=2.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.01051
.param par_k=0.00517
.param par_l=3e-7
.param par_w=-4e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b pplus_u_m2 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b pplus_u_m2 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b pmos_6p0 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='0' sb='0' sd='0' delvto='mis_vth*sw_stat_mismatch'
.ends
.model pmos_6p0.0 pmos a0=0.84 a1=0 a2=1 acde=0.7 acnqsmod=0 agidl=1.1e-15 ags=0.059 alpha0=9.6e-7 alpha1=51.5 at=-2.18e4 b0=2.625e-8 b1=0 beta0=50.8 bgidl=1.578e5 binunit=1 bvd=10.5 bvs=10.5 capmod=2 cdsc=2.4e-4 cdscb=0 cdscd=0 cgbo=1e-13 cgdl='5.25e-11*pmos_6p0_dcgdo' cgdo='7.71e-11*pmos_6p0_dcgdo' cgsl='5.25e-11*pmos_6p0_dcgso' cgso='7.71e-11*pmos_6p0_dcgso' cit=0 cjd=0.000912 cjs=0.000912 cjswd=1.4649e-010 cjswgd=3.3229e-010 cjswgs=3.3229e-010 cjsws=1.4649e-010 ckappad=0.6 ckappas=0.6 delta=0.01 diomod=1 dlc=7.4e-9 drout=0.56 dsub=0.4824 dvt0=1 dvt0w=0 dvt1=1 dvt1w=5.3e6 dvt2=0 dvt2w=-0.032 dvtp0=0 dvtp1=0.3 dwb=-3e-9 dwg=-6.6e-9 ef=1.1 egidl=1.19653e-2 epsrox=3.9 eta0=0.08 etab=-0.09408 fnoimod=1 fprout=0 geomod=1 igbmod=0 igcmod=0 ijthdfwd=0.1 ijthdrev=0.1 ijthsfwd=0.1 ijthsrev=0.1 jsd=2.0867e-007 jss=2.0867e-007 jswd=1.6088e-013 jswgd=0 jswgs=0 jsws=1.6088e-013 k1=0.9588 k2=8.936e-3 k3=-0.75 k3b=1.2104 keta=-8.6016e-5 kt1=-0.3828 kt1l=-3.158e-8 kt2=-0.09064 lambda=0 lc=0 level=54 lint=6.7e-8 ll=-5.4e-15 lln=1 lmax=50.01e-6 lmin=0.5e-6 lpe0=-4.4e-8 lpeb=-5.96e-8 lphin=0.1408 lua1=-6.554813e-10 lub1=1.939773e-19 luc1=-1.067674e-10 luc=8.691408e-11 lute=-0.152467 lw=0 lwl=-4.76e-21 lwn=1 minv=0 mjd=0.32713 mjs=0.32713 mjswd=0.056777 mjswgd=0.50996 mjswgs=0.50996 mjsws=0.056777 mobmod=0 moin=15 ndep=1.7e17 nfactor=1 ngate=3.6e19 njd=1 njs=1 noff=1 noia='pmos_6p0_noia' noib='pmos_6p0_noib' noic='pmos_6p0_noic' nsd=6e16 pagidl=6.27545e-16 paramchk=1 pat=-6.1e3 pbd=0.76836 pbeta0=0.14 pbs=0.76836 pbswd=0.5 pbswgd=1.2295 pbswgs=1.2295 pbsws=0.5 pclm=0.42 pdiblc1=0.14 pdiblc2=1e-5 pdiblcb=0 pdits=0.01 pditsd=0 pditsl=0 permod=1 petab=-0.012128 phin=0 pkt1=2.2e-3 ppclm=0.071 pprwb=-0.052 prdsw=-120 prt=454 prwb=0.569552 prwg=0.0432 pscbe1=5.088e8 pscbe2=1e-8 pua1=-3.823641e-10 pub1=7.291324e-19 puc1=1.8536e-11 puc=-1.501336e-11 pvag=1.5 pvth0='7.6e-3+8.47e-3*pmos_6p0_dvth0' rbodymod=0 rdsmod=0 rdsw=1.426e3 rdswmin=100 rsh=7 rshg=0.1 tcj=0.001 tcjsw=0.00071888 tcjswg=0.0009411 tempmod=0 tnoimod=0 tnom=25 toxe='1.56e-8+pmos_6p0_dtox' tpb=0.0019314 tpbsw=0.0017642 tpbswg=0.0016588 trnqsmod=0 u0=0.0151 ua1=1.41e-9 ua=1.78e-9 ub1=-4.31e-18 ub=4.88e-19 uc1=1.147552e-10 uc=-2.7435e-11 ute=-1.2 version=4.5 vfb=-1 voff=-0.1284 voffcv=0 voffl=2.19e-8 vsat=8.55e4 vth0='-0.8978+pmos_6p0_dvth0' vtl=2e5 w0=3.1e-7 wbeta0=0.22 wint=4.9e-8 wketa=2.772e-3 wl=0 wln=1 wmax=100.01e-6 wmin=0.3e-6 wr=1 wrdsw=213.9 wua1=-1.2e-10 wute=-0.07 ww=-1.37e-14 wwl=3.04e-22 wwn=1 xj=1.5e-7 xjbvd=1 xjbvs=1 xl='0+pmos_6p0_dxl' xn=3 xpart=1 xtid=3 xtis=3 xw='0+pmos_6p0_dxw'
.subckt pplus_u_m2 1 2 3 r_length='lr' r_width='wr' dtemp=0 par=1 r_rsh0='rsh_pplus_u_m' r_dw=2.75e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.375e-3 r_tc2=1e-6 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model pn_junction d cj=0.00094344 level=2
d1 1 3 pn_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends pplus_u_m2
.endl pmos_6p0_t

.lib dio
.model np_3p3 d cj='0.00096797*cja' eg=1.17 ibv=0.001 is='2.2959e-007*jsa' n=1.01 rs='2e-010*rsa' bv=11.0 xti=3 tnom=25 ikf=300000 level=2
.model pn_3p3 d cj='0.00094344*cja' eg=1.17 ibv=0.001 is='1.653e-007*jsa' n=1 rs='2e-010*rsa' bv=10.5 xti=3 level=2
.model np_6p0 d cj='0.00095*cja' eg=1.11 ibv=0.001 is='6.88e-007*jsa' n=1.0541 rs='2e-010*rsa' bv=11 xti=5 level=2
.model pn_6p0 d bv=10.5 cj='0.000912*cja' eg=1.17 is='2.0867e-007*jsa' n=1.0058 rs='2.0e-010*rsa' xti=3 level=2
.model nwp_3p3 d cj='0.00014917*cja' eg=1.18 ibv=0.001 is='1.5654e-006*jsa' n=1.01 rs='2e-010*rsa' bv=14 xti=3 level=2
.model nwp_6p0 d bv=14 cj='0.00014914*cja' eg=1.1763 is='1.6119e-006*jsa' n=1 rs='2e-010*rsa' xti=3 level=2
.model dnwpw d cj='0.00032124*cja' eg=1.17 ibv=0.001 is='5.2139e-007*jsa' n=0.98 rs='2e-010*rsa' bv=14.732 xti=3 level=2
.model dnwps d cj='0.00022998*cja' eg=1.17 ibv=0.001 is='2e-006*jsa' n=0.99335 rs='2e-010*rsa' bv=30.48 xti=3 level=2
.model sc_diode d cj='0.00176*cja_sc' eg=0.61 ibv=9.92e-005 js='8.16*10**jsa_sc' n=1.0553 rs='2.768e-009*rs_sc' bv='17+vba_sc' xti=3 level=2
.endl dio

.lib res
.subckt nplus_u 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_nplus_u*(1+(mc_rsh_nplus_u/(rsh_nplus_u))*res_mc_skew*sw_stat_global)' r_dw='-5e-8*(1+mc_dw_nplus_u*res_mc_skew*sw_stat_global)' r_dl=2e-11 r_vc1=0 r_vc2=0 r_tc1=1.36e-3 r_tc2=6.5e-7 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)' par_r=0.012608 par_sqrtarea='sqrt(par*(r_l)*(r_w))' var_r='0.7071*par_r*1e-06/par_sqrtarea' mis_r='agauss(0,var_r,1)'
.model nplus_u_t r rsh='18.5+mc_rt_nplus_u*res_mc_skew*sw_stat_global' tc1=8.5e-4 tc2=1.75e-6 level=1
.model np_3p3 d cj=0.00096797 level=2
rt1 1 11 nplus_u_t l='s*1u' w='r_w'
d1 3 1 np_3p3 area='r_w*r_l/2'
rb 11 21 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)*(1+mis_r*sw_stat_mismatch)'
rt2 21 2 nplus_u_t l='s*1u' w='r_w'
d2 3 2 np_3p3 area='r_w*r_l/2'
.ends nplus_u
.subckt pplus_u 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_pplus_u*(1+mc_rsh_pplus_u/(rsh_pplus_u)*res_mc_skew*sw_stat_global)' r_dw='2.75e-8*(1+mc_dw_pplus_u*res_mc_skew*sw_stat_global)' r_dl=5.0e-11 r_vc1=0 r_vc2=0 r_tc1=1.375e-3 r_tc2=1e-6 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)' par_r=0.0126 par_sqrtarea='sqrt(par*(r_l)*(r_w))' var_r='0.7071*par_r*1e-06/par_sqrtarea' mis_r='agauss(0,var_r,1)'
.model pplus_u_t r rsh='50+mc_rt_pplus_u*res_mc_skew*sw_stat_global' tc1=-1.528e-3 tc2=0.7e-6 level=1
.model pn_3p3 d cj=0.00094344 level=2
rt1 1 11 pplus_u_t l='s*1u' w='r_w'
d1 1 3 pn_3p3 area='r_w*r_l/2'
rb 11 21 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)*(1+mis_r*sw_stat_mismatch)'
rt2 21 2 pplus_u_t l='s*1u' w='r_w'
d2 2 3 pn_3p3 area='r_w*r_l/2'
.ends pplus_u
.subckt nplus_s 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_nplus_s*(1+mc_rsh_nplus_s/(rsh_nplus_s)*res_mc_skew*sw_stat_global)' r_dw='-1.25e-8*(1+mc_dw_nplus_s*res_mc_skew*sw_stat_global)' r_dl=3.5e-11 r_vc1=0 r_vc2=0 r_tc1=3.3e-3 r_tc2=3e-7 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model nplus_s_t r rsh=6 tc1=1.43e-3 tc2=-0.27e-6 level=1
.model np_3p3 d cj=0.00096797 level=2
rt1 1 11 nplus_s_t l='s*1u' w='r_w'
d1 3 1 np_3p3 area='r_w*r_l/2'
rb 11 21 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)'
rt2 21 2 nplus_s_t l='s*1u' w='r_w'
d2 3 2 np_3p3 area='r_w*r_l/2'
.ends nplus_s
.subckt pplus_s 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_pplus_s*(1+mc_rsh_pplus_s/(rsh_pplus_s)*res_mc_skew*sw_stat_global)' r_dw='-5e-8*(1+mc_dw_pplus_s*res_mc_skew*sw_stat_global)' r_dl=3.5e-11 r_vc1=0 r_vc2=0 r_tc1=3.375e-3 r_tc2=0.45e-6 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model pplus_s_t r rsh=6.5 tc1=1.565e-3 tc2=-0.028e-6 level=1
.model pn_3p3 d cj=0.00094344 level=2
rt1 1 11 pplus_s_t l='s*1u' w='r_w'
d1 1 3 pn_3p3 area='r_w*r_l/2'
rb 11 21 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)'
rt2 21 2 pplus_s_t l='s*1u' w='r_w'
d2 2 3 pn_3p3 area='r_w*r_l/2'
.ends pplus_s
.subckt nwell 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_nwell' r_dw=2.22e-7 r_dl=1.02e-8 r_vc1=0 r_vc2=0 r_tc1=2.285e-3 r_tc2=9.78e-6 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model nwell_t r rsh=250 tc1=1.72e-3 tc2=9.34e-6 level=1
.model nwp d cj=0.00014917 level=2
rt1 1 11 nwell_t l='s*1u' w='r_w'
d1 3 1 nwp area='r_w*r_l/2'
rb 11 21 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)'
rt2 21 2 nwell_t l='s*1u' w='r_w'
d2 3 2 nwp area='r_w*r_l/2'
.ends nwell
.subckt npolyf_u 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_npolyf_u*(1+mc_rsh_npolyf_u/(rsh_npolyf_u)*res_mc_skew*sw_stat_global)' r_dw='0.0265e-6*(1+mc_dw_npolyf_u*res_mc_skew*sw_stat_global)' r_dl=8.48e-11 r_vc1=0 r_vc2=0 r_tc1=-1.4e-3 r_tc2=2.2e-6 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)' par_r=0.05808 par_sqrtarea='sqrt(par*(r_l)*(r_w))' var_r='0.7071*par_r*1e-06/par_sqrtarea' mis_r='agauss(0,var_r,1)'
.model npolyf_u_body r level=1
.model npolyf_u_t r rsh='40+mc_rt_npolyf_u*res_mc_skew*sw_stat_global' tc1=-0.735e-3 tc2=-1.7e-6 level=1
.model fox_sub c cj=8.85e-05
rt1 1 11 npolyf_u_t l='s*1u' w='r_w'
c1 1 3 fox_sub l='r_l/2' w='r_w'
rb 11 21 npolyf_u_body r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)*(1+mis_r*sw_stat_mismatch)' l='r_l' w='r_w'
rt2 21 2 npolyf_u_t l='s*1u' w='r_w'
c2 2 3 fox_sub l='r_l/2' w='r_w'
.ends npolyf_u
.subckt ppolyf_u 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_ppolyf_u*(1+mc_rsh_ppolyf_u/(rsh_ppolyf_u)*res_mc_skew*sw_stat_global)' r_dw='2.55e-8*(1+mc_dw_ppolyf_u*res_mc_skew*sw_stat_global)' r_dl=2e-11 r_vc1=0 r_vc2=0 r_tc1=-0.9e-4 r_tc2=7e-7 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)' par_r=0.021 par_sqrtarea='sqrt(par*(r_l)*(r_w))' var_r='0.7071*par_r*1e-06/par_sqrtarea' mis_r='agauss(0,var_r,1)'
.model ppolyf_u_body r level=1
.model ppolyf_u_t r rsh='60+mc_rt_ppolyf_u*res_mc_skew*sw_stat_global' tc1=-1.47e-3 tc2=0.82e-6 level=1
.model fox_sub c cj=8.85e-05
rt1 1 11 ppolyf_u_t l='s*1u' w='r_w'
c1 1 3 fox_sub l='r_l/2' w='r_w'
rb 11 21 ppolyf_u_body r='(r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n))*(1+mis_r*sw_stat_mismatch)' l='r_l' w='r_w'
rt2 21 2 ppolyf_u_t l='s*1u' w='r_w'
c2 2 3 fox_sub l='r_l/2' w='r_w'
.ends ppolyf_u
.subckt npolyf_s 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_npolyf_s*(1+mc_rsh_npolyf_s/(rsh_npolyf_s)*res_mc_skew*sw_stat_global)' r_dw='6.5e-9*(1+mc_dw_npolyf_s*res_mc_skew*sw_stat_global)' r_dl=1.5e-11 r_vc1=0 r_vc2=0 r_tc1=3.26e-3 r_tc2=0.25e-6 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model npolyf_s_body r level=1
.model npolyf_s_t r rsh=5.5 tc1=1.28e-3 tc2=-0.5e-6 level=1
.model fox_sub c cj=8.85e-05
rt1 1 11 npolyf_s_t l='s*1u' w='r_w'
c1 1 3 fox_sub l='r_l/2' w='r_w'
rb 11 21 npolyf_s_body r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)' l='r_l' w='r_w'
rt2 21 2 npolyf_s_t l='s*1u' w='r_w'
c2 2 3 fox_sub l='r_l/2' w='r_w'
.ends npolyf_s
.subckt ppolyf_s 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_ppolyf_s*(1+mc_rsh_ppolyf_s/(rsh_ppolyf_s)*res_mc_skew*sw_stat_global)' r_dw='7.5e-9*(1+mc_dw_ppolyf_s*res_mc_skew*sw_stat_global)' r_dl=1.5e-10 r_vc1=0 r_vc2=0 r_tc1=3.245e-3 r_tc2=3.6e-7 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model ppolyf_s_body r level=1
.model ppolyf_s_t r rsh=5 tc1=1.254e-3 tc2=-0.27e-6 level=1
.model fox_sub c cj=8.85e-05
rt1 1 11 ppolyf_s_t l='s*1u' w='r_w'
c1 1 3 fox_sub l='r_l/2' w='r_w'
rb 11 21 ppolyf_s_body r='(r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n))' l='r_l' w='r_w'
rt2 21 2 ppolyf_s_t l='s*1u' w='r_w'
c2 2 3 fox_sub l='r_l/2' w='r_w'
.ends ppolyf_s
.subckt ppolyf_u_1k 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1
.param r_rsh0='rsh_ppolyf_u_1k*(1+mc_rsh_ppolyf_u_1k/(rsh_ppolyf_u_1k)*res_mc_skew*sw_stat_global)'
.param r_dw='0.0148e-6*(1+mc_dw_ppolyf_u_1k*res_mc_skew*sw_stat_global)'
.param r_dl=3.85e-11
.param r_vc1=0
.param r_vc2=0
.param r_tc1=-9.39e-4
.param r_tc2=2.51e-6
.param r_tnom=25
.param r_l='s*(r_length-2*r_dl)'
.param r_w='r_width-2*r_dw'
.param r_n='r_l/r_w'
.param r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model ppolyf_u_1k_body r level=1
.model ppolyf_u_1k_t r rsh='85.45+mc_rt_ppolyf_u_1k*res_mc_skew*sw_stat_global' tc1=-7.92e-3 tc2=4.25e-5 level=1
.model fox_sub c cj=8.85e-05
rt1 1 11 ppolyf_u_1k_t l='s*1u' w='r_w'
c1 1 3 fox_sub l='r_l/2' w='r_w'
rb 11 21 ppolyf_u_1k_body r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)' l='r_l' w='r_w'
rt2 21 2 ppolyf_u_1k_t l='s*1u' w='r_w'
c2 2 3 fox_sub l='r_l/2' w='r_w'
.ends ppolyf_u_1k
.subckt ppolyf_u_2k 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1
.param r_rsh0='rsh_ppolyf_u_2k*(1+mc_rsh_ppolyf_u_2k/(rsh_ppolyf_u_2k)*res_mc_skew*sw_stat_global)'
.param r_dw='0.02256e-6*(1+mc_dw_ppolyf_u_2k*res_mc_skew*sw_stat_global)'
.param r_dl=-0.0932e-6
.param r_vc1=0
.param r_vc2=0
.param r_tc1=-0.001669823
.param r_tc2=3.74326e-06
.param r_tnom=25
.param r_l='s*(r_length-2*r_dl)'
.param r_w='r_width-2*r_dw'
.param r_n='r_l/r_w'
.param r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model ppolyf_u_2k_body r level=1
.model ppolyf_u_2k_t r rsh='33.16+mc_rt_ppolyf_u_2k*res_mc_skew*sw_stat_global' tc1=-0.003763316 tc2=9.81166e-06 level=1
.model fox_sub c cj=8.85e-05
rt1 1 11 ppolyf_u_2k_t l='s*1u' w='r_w'
c1 1 3 fox_sub l='r_l/2' w='r_w'
rb 11 21 ppolyf_u_2k_body r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)' l='r_l' w='r_w'
rt2 21 2 ppolyf_u_2k_t l='s*1u' w='r_w'
c2 2 3 fox_sub l='r_l/2' w='r_w'
.ends ppolyf_u_2k
.subckt ppolyf_u_1k_6p0 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1
.param r_rsh0='rsh_ppolyf_u_1k_6p0*(1+mc_rsh_ppolyf_u_1k_6p0/(rsh_ppolyf_u_1k_6p0)*res_mc_skew*sw_stat_global)'
.param r_dw='0.0148e-6*(1+mc_dw_ppolyf_u_1k_6p0*res_mc_skew*sw_stat_global)'
.param r_dl=3.85e-11
.param r_vc1=0
.param r_vc2=0
.param r_tc1=-9.39e-4
.param r_tc2=2.51e-6
.param r_tnom=25
.param r_l='s*(r_length-2*r_dl)'
.param r_w='r_width-2*r_dw'
.param r_n='r_l/r_w'
.param r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model ppolyf_u_1k_body r level=1
.model ppolyf_u_1k_t r rsh='85.45+mc_rt_ppolyf_u_1k_6p0*res_mc_skew*sw_stat_global' tc1=-7.92e-3 tc2=4.25e-5 level=1
.model fox_sub c cj=8.85e-05
rt1 1 11 ppolyf_u_1k_t l='s*1u' w='r_w'
c1 1 3 fox_sub l='r_l/2' w='r_w'
rb 11 21 ppolyf_u_1k_body r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)' l='r_l' w='r_w'
rt2 21 2 ppolyf_u_1k_t l='s*1u' w='r_w'
c2 2 3 fox_sub l='r_l/2' w='r_w'
.ends ppolyf_u_1k_6p0
.subckt ppolyf_u_2k_6p0 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1
.param r_rsh0='rsh_ppolyf_u_2k_6p0+mc_rsh_ppolyf_u_2k_6p0*res_mc_skew*sw_stat_global'
.param r_dw='0.02256e-6*(1+mc_dw_ppolyf_u_2k_6p0*res_mc_skew*sw_stat_global)'
.param r_dl=-0.0932e-6
.param r_vc1=0
.param r_vc2=0
.param r_tc1=-0.001669823
.param r_tc2=3.74326e-06
.param r_tnom=25
.param r_l='s*(r_length-2*r_dl)'
.param r_w='r_width-2*r_dw'
.param r_n='r_l/r_w'
.param r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model ppolyf_u_2k_body r level=1
.model ppolyf_u_2k_t r rsh='33.16+mc_rt_ppolyf_u_2k_6p0*res_mc_skew*sw_stat_global' tc1=-0.003763316 tc2=9.81166e-06 level=1
.model fox_sub c cj=8.85e-05
rt1 1 11 ppolyf_u_2k_t l='s*1u' w='r_w'
c1 1 3 fox_sub l='r_l/2' w='r_w'
rb 11 21 ppolyf_u_2k_body r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)' l='r_l' w='r_w'
rt2 21 2 ppolyf_u_2k_t l='s*1u' w='r_w'
c2 2 3 fox_sub l='r_l/2' w='r_w'
.ends ppolyf_u_2k_6p0
.subckt ppolyf_u_3k 1 2 3 r_length='l' r_width='w' dtemp=0 par=1 s=1
.param r_rsh0='rsh_ppolyf_u_3k*(1+mc_rsh_ppolyf_u_3k/(rsh_ppolyf_u_3k)*res_mc_skew*sw_stat_global)'
.param r_dw='0.02256e-6*(1+mc_dw_ppolyf_u_3k*res_mc_skew*sw_stat_global)'
.param r_dl=-0.0932e-6
.param r_vc1=0
.param r_vc2=0
.param r_tc1=-0.001669823
.param r_tc2=3.74326e-06
.param r_tnom=25
.param r_l='s*(r_length-2*r_dl)'
.param r_w='r_width-2*r_dw'
.param r_n='r_l/r_w'
.param r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model ppolyf_u_3k_body r level=1
.model ppolyf_u_3k_t r rsh='33.16+mc_rt_ppolyf_u_3k*res_mc_skew*sw_stat_global' tc1=-0.003763316 tc2=9.81166e-06 level=1
.model fox_sub c cj=8.85e-05
rt1 1 11 ppolyf_u_3k_t l='s*1u' w='r_w'
c1 1 3 fox_sub l='r_l/2' w='r_w'
rb 11 21 ppolyf_u_3k_body r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(11,21))/r_n+r_vc2*abs(v(11,21))*abs(v(11,21))/r_n/r_n)' l='r_l' w='r_w'
rt2 21 2 ppolyf_u_3k_t l='s*1u' w='r_w'
c2 2 3 fox_sub l='r_l/2' w='r_w'
.ends ppolyf_u_3k
.subckt rm1 1 2 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_rm1' r_dw=0 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=3.33e-3 r_tc2=0 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends rm1
.subckt rm2 1 2 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_rm2' r_dw=0 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=3.33e-3 r_tc2=0 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends rm2
.subckt rm3 1 2 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_rm3' r_dw=0 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=3.33e-3 r_tc2=0 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends rm3
.subckt tm6k 1 2 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_tm6k' r_dw=0 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=3.5e-3 r_tc2=0 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends tm6k
.subckt tm9k 1 2 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_tm9k' r_dw=0 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=3.7e-3 r_tc2=0 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends tm9k
.subckt tm11k 1 2 r_length='l' r_width='w' dtemp=0 par=1 s=1 r_rsh0='rsh_tm11k' r_dw=0 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=3.7e-3 r_tc2=0 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends tm11k
.subckt tm30k 1 2 r_length='l' r_width='w' par=1 s=1 dtemp=0 r_rsh0='rsh_tm30k' r_dw=0 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=3.86e-3 r_tc2=1.51e-6 r_tnom=25 r_l='s*(r_length-2*r_dl)' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends tm30k
.endl res

.lib mim_cap
.subckt mim_1p5ff 1 2 c_length='l' c_width='w' dtemp=0 par=1
.param c_cox='1.47e-3*mim_corner_1p5ff'
.param c_capsw='3.79e-10*mim_corner_1p5ff'
.param c_tnom=25
.param c_tc1=4.0604e-05
.param c_tc2=-6.90e-08
.param c_vcr1=-4.5152e-05
.param c_vcr2=9.748e-06
.param c_area='c_length*c_width'
.param c_peri='2*(c_length+c_width)'
.param c_c0='(c_cox*c_area+c_capsw*c_peri)*(1+c_tc1*(temp+dtemp-c_tnom)+c_tc2*(temp+dtemp-c_tnom)*(temp+dtemp-c_tnom))'
c_cap 1 2 c='c_c0*(1+c_vcr1*v(1,2)+c_vcr2*v(1,2)*v(1,2))*(1+mc_c_cox_1p5ff)'
.ends mim_1p5ff
.subckt mim_1p0ff 1 2 c_length='l' c_width='w' dtemp=0 par=1
.param c_cox='0.987e-3*mim_corner_1p0ff'
.param c_capsw='3.3e-10*mim_corner_1p0ff'
.param c_tnom=25
.param c_tc1=1.302e-5
.param c_tc2=-4.93e-9
.param c_vcr1=6.079e-6
.param c_vcr2=1.268e-6
.param c_area='c_length*c_width'
.param c_peri='2*(c_length+c_width)'
.param c_c0='(c_cox*c_area+c_capsw*c_peri)*(1+c_tc1*(temp+dtemp-c_tnom)+c_tc2*(temp+dtemp-c_tnom)*(temp+dtemp-c_tnom))'
c_cap 1 2 c='c_c0*(1+c_vcr1*v(1,2)+c_vcr2*v(1,2)*v(1,2))*(1+mc_c_cox_1p0ff)'
.ends mim_1p0ff
.subckt mim_2p0ff 1 2 c_length='l' c_width='w' dtemp=0 par=1
.param gleak='9.51e-10/5*10000'
.param c_cox='1.99e-3*mim_corner_2p0ff'
.param c_capsw='2.383e-10*mim_corner_2p0ff'
.param c_vcr1='0+(c_width>5u||c_length>5u)*8.742e-6+(c_width<=5u||c_length<=5u)*(-81e-6)'
.param c_vcr2='0+(c_width>5u||c_length>5u)*9.188e-6+(c_width<=5u||c_length<=5u)*(16.7e-6)'
.param c_tnom=25
.param c_tc1=1.46e-5
.param c_tc2=-5.55e-8
.param c_area='c_length*c_width'
.param c_peri='2*(c_length+c_width)'
.param c_c0='(c_cox*c_area+c_capsw*c_peri)*(1+c_tc1*(temp+dtemp-c_tnom)+c_tc2*(temp+dtemp-c_tnom)*(temp+dtemp-c_tnom))'
c_cap 1 2 c='c_c0*(1+c_vcr1*v(1,2)+c_vcr2*v(1,2)*v(1,2))*(1+mc_c_cox_2p0ff)'
r_leak 1 2 r='1/(gleak*c_area)' tc1='c_tc1' tc2='c_tc2'
.ends mim_2p0ff
.endl mim_cap

.lib moscap
.subckt nmoscap_3p3 1 2 c_length='l' c_width='w' dtemp=0
.param cvar1=0.002003
.param cvar2=0.00198
.param cvar3=6.25
.param cvar4=-3.9375
c_moscap 1 2 c='nmoscap_3p3_corner*l*w*(cvar1+cvar2*tanh(cvar3*v(1,2)+cvar4))'
.ends nmoscap_3p3
.subckt pmoscap_3p3 1 2 c_length='l' c_width='w' dtemp=0
.param cvar1=0.001998
.param cvar2=0.00196
.param cvar3=-6.25
.param cvar4=-4.9375
c_moscap 1 2 c='pmoscap_3p3_corner*l*w*(cvar1+cvar2*tanh(cvar3*v(1,2)+cvar4))'
.ends pmoscap_3p3
.subckt nmoscap_6p0 1 2 c_length='l' c_width='w' dtemp=0
.param cvar1=0.001107
.param cvar2=0.00107
.param cvar3=6.25
.param cvar4=-4.1875
c_moscap 1 2 c='nmoscap_6p0_corner*l*w*(cvar1+cvar2*tanh(cvar3*v(1,2)+cvar4))'
.ends nmoscap_6p0
.subckt pmoscap_6p0 1 2 c_length='l' c_width='w' dtemp=0
.param cvar1=0.001107
.param cvar2=0.00107
.param cvar3=-6.25
.param cvar4=-5.75
c_moscap 1 2 c='pmoscap_6p0_corner*l*w*(cvar1+cvar2*tanh(cvar3*v(1,2)+cvar4))'
.ends pmoscap_6p0
.subckt nmoscap_3p3_b 1 2 c_length='l' c_width='w' dtemp=0
.param cvar1=0.002458
.param cvar2=0.001533
.param cvar3=1.515152
.param cvar4=0.560606
c_moscap 1 2 c='nmoscap_3p3_b_corner*l*w*(cvar1+cvar2*tanh(cvar3*v(1,2)+cvar4))'
.ends nmoscap_3p3_b
.subckt pmoscap_3p3_b 1 2 c_length='l' c_width='w' dtemp=0
.param cvar1=0.002435
.param cvar2=0.00154
.param cvar3=-1.66667
.param cvar4=0.65
c_moscap 1 2 c='pmoscap_3p3_b_corner*l*w*(cvar1+cvar2*tanh(cvar3*v(1,2)+cvar4))'
.ends pmoscap_3p3_b
.subckt nmoscap_6p0_b 1 2 c_length='l' c_width='w' dtemp=0
.param cvar1=0.001293
.param cvar2=0.000863
.param cvar3=1.052632
.param cvar4=0.736842
c_moscap 1 2 c='nmoscap_6p0_b_corner*l*w*(cvar1+cvar2*tanh(cvar3*v(1,2)+cvar4))'
.ends nmoscap_6p0_b
.subckt pmoscap_6p0_b 1 2 c_length='l' c_width='w' dtemp=0
.param cvar1=0.001325
.param cvar2=0.000865
.param cvar3=-1.42857
.param cvar4=0.642857
c_moscap 1 2 c='pmoscap_6p0_b_corner*l*w*(cvar1+cvar2*tanh(cvar3*v(1,2)+cvar4))'
.ends pmoscap_6p0_b
.endl moscap

.lib nmos_3p3_stat
.subckt nmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.007148
.param par_k=0.007008
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b nplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b nplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b nmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model nmos_3p3.0 nmos a0=0.11197377 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.32403844 alpha0=2.652013e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=19.905584 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0036363636 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95938091 k2=0.054714558 k3=0 k3b=0 keta=-0.14896036 kt1=-0.45934558 kt1l=0 kt2=-0.024730519 ku0=0 kvsat=0 kvth0=0 la0=-3.1454545e-009 lags=-1.5116364e-008 lalpha0=-3.0506364e-013 lbeta0=1.2863636e-007 ldelta=3.1818182e-009 level=54 lint=0 lk1=-9.9985454e-008 lk2=-4.1647636e-008 lketa=3.8830182e-008 lkt1=4.2126364e-008 lkt2=1.2545455e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-4.729e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.6525455e-009 lua=7.0220545e-016 lub1=2.8745455e-025 lub=-7.9058636e-025 luc1=-3.8181818e-018 luc=-6.1360545e-017 lute=9.0909091e-008 lvoff=3.9354545e-009 lvsat=-0.0027272727 lvth0=-3.8715455e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.7450182e-015 pags=-1.2213818e-014 palpha0=-1.3658182e-020 paramchk=1 pbeta0=8.7272727e-016 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.3741 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=5.388e-015 pketa=-2.4261818e-015 pkt1=-8.6530909e-015 pkt2=-2.9672727e-016 ppclm=8.5658182e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-6.5127273e-016 pua=-1.4149745e-022 pub1=-5.7490909e-032 pub=9.2644364e-032 puc1=1.8327273e-024 puc=5.4467782e-024 pute=-4.3636364e-014 pvag=0 pvoff=-1.4858182e-015 pvsat=1.3090909e-009 pvth0=4.3636364e-016 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.023671338 ua1=1.675e-009 ua=-1.1554452e-009 ub1=-4.1945234e-018 ub=3.3771156e-018 uc1=-4.2363636e-011 uc=2.2660166e-010 ute=-1.5675325 vbm=-3 version=4.5 vfbcv=-1 voff=-0.1262652 voffcv=0.005 voffl=0 vsat=92454.546 vth0='nmos_3p3_vth0_0' w0=5e-007 wa0=-6.2322078e-009 wags=4.7930493e-008 walpha0=4.8779221e-014 wbeta0=1.3848312e-007 wint=1e-008 wk2=-1.9242857e-008 wketa=8.1643636e-009 wkt1=3.2086753e-008 wkt2=1.0597403e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.1028364e-008 wr=1 wtvoff=0 wu0=4.6066597e-009 wua=2.7073777e-016 wub1=3.3492467e-025 wub=-4.093733e-025 wuc1=-6.5454545e-018 wuc=-3.2577351e-017 wute=1.0441558e-007 wvoff=5.3064935e-009 wvsat=-0.00021818182 wvth0=-1.430587e-008 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.1 nmos a0=1.0861147 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.47870122 alpha0=6.5720816e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=22.625306 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0014285714 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.74639857 k2=0.0237458 k3=0 k3b=0 keta=-0.028417143 kt1=-0.33916633 kt1l=0 kt2=-0.020311225 ku0=0 kvsat=0 kvth0=0 la0=-4.9021592e-007 lags=-9.2447755e-008 lalpha0=-2.265098e-012 lbeta0=-1.2312245e-006 ldelta=4.2857143e-009 level=54 lint=0 lk1=6.5057143e-009 lk2=-2.6163257e-008 lketa=-2.1441429e-008 lkt1=-1.7963265e-008 lkt2=-9.5510204e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=9.8313061e-008 lpdiblc2=9.06e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.6503673e-009 lua=7.7258204e-016 lub1=-4.0760816e-025 lub=-6.4387347e-025 luc1=5.1428571e-018 luc=9.6333061e-018 lvoff=-2.8273469e-009 lvsat=0.0017142857 lvth0=-2.3433061e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.4627526e-014 pags=-9.9007347e-015 palpha0=1.8396735e-020 paramchk=1 pbeta0=2.4538775e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.082893878 pdiblc1=0.39 pdiblc2=0.001359 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=-2.7269486e-015 pketa=5.3691429e-015 pkt1=8.6223674e-015 pkt2=2.5273469e-016 ppclm=-2.8711837e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.2234122e-015 pua=-2.976098e-023 pub1=8.1521633e-032 pub=-9.8501878e-032 puc1=-2.4685714e-024 puc=-1.1961815e-023 pvag=0 pvoff=3.2032653e-016 pvsat=2.0571429e-009 pvth0=-5.642449e-016 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.029675694 ua1=1.675e-009 ua=-1.2961984e-009 ub1=-2.804398e-018 ub=3.0836898e-018 uc1=-6.0285714e-011 uc=8.4613959e-011 ute=-1.3857143 vbm=-3 version=4.5 vfbcv=-1 voff=-0.11273959 voffcv=0.005 voffl=0 vsat=83571.429 vth0='nmos_3p3_vth0_1' w0=5e-007 wa0=-5.1997224e-008 wags=4.3304327e-008 walpha0=-1.5330612e-014 wbeta0=-3.5054694e-007 wint=1e-008 wk2=-3.01296e-009 wketa=-7.4262857e-009 wkt1=-2.4641633e-009 wkt2=-3.9183673e-011 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=4.3902367e-008 wr=1 wtvoff=0 wu0=8.572898e-010 wua=4.7264816e-017 wub1=5.6899592e-026 wub=-2.7080816e-026 wuc1=2.0571429e-018 wuc=2.2398367e-018 wute=1.7142857e-008 wvoff=1.6942041e-009 wvsat=-0.0017142857 wvth0=-1.2304653e-008 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.2 nmos a0=1.224418 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.25784649 alpha0=7.5243347e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.210162 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027272727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79593364 k2=0.0056393844 k3=0 k3b=0 keta=-0.019651071 kt1=-0.32898149 kt1l=0 kt2=-0.021107143 ku0=0 kvsat=0 kvth0=0 la0=-6.5617987e-007 lags=1.7257792e-007 lalpha0=-8.4670617e-011 lbeta0=-3.133052e-006 ldelta=2.7272727e-009 level=54 lint=0 lk1=-5.2936364e-008 lk2=-4.4355584e-009 lketa=-3.1960714e-008 lkt1=-3.0185065e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=-2.9236364e-008 lpdiblc2=1.7686364e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.6755195e-009 lua=1.9570909e-016 lub1=-7.5296104e-025 lub=-2.347987e-025 luc=-6.9921429e-018 lvoff=1.3461039e-008 lvth0=-3.224026e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-4.2919481e-014 pags=4.5191688e-014 palpha0=-9.043013e-018 paramchk=1 pbeta0=-3.1184416e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.18918506 pdiblc1=0.39 pdiblc2=0.00064013636 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=2.6091117e-015 pketa=-2.7504935e-015 pkt1=1.4488831e-014 ppclm=4.7225454e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.447013e-015 pua=1.9701818e-023 pub1=1.231013e-031 pub=-1.1174026e-031 puc=1.4030649e-024 pvag=0 pvoff=-1.4493507e-016 pvth0=-3.6888312e-015 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032447266 ua1=1.675e-009 ua=-8.1547091e-010 ub1=-2.5166039e-018 ub=2.7427942e-018 uc1=-5.6e-011 uc=9.84685e-011 ute=-1.3857143 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12631325 voffcv=0.005 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_2' w0=5e-007 wa0=4.291948e-009 wags=-2.606026e-009 walpha0=7.5358442e-012 wbeta0=1.1381299e-007 wint=1e-008 wk2=-7.4596769e-009 wketa=-6.5992208e-010 wkt1=-7.3528831e-009 wkt2=1.7142857e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.1551688e-009 wr=1 wtvoff=0 wu0=6.7095584e-010 wua=6.0458182e-018 wub1=2.224987e-026 wub=-1.6048831e-026 wuc=-8.8975636e-018 wute=1.7142857e-008 wvoff=2.0819221e-009 wvth0=-9.7008312e-009 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.3 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.27510429 alpha0=6.6776286e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.896857 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=0.0051958286 k3=0 k3b=0 keta=-0.022847143 kt1=-0.332 kt1l=0 kt2=-0.021107143 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.18626143 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.032279714 ua1=1.675e-009 ua=-7.959e-010 ub1=-2.5919e-018 ub=2.7193143e-018 uc1=-5.6e-011 uc=9.7769286e-011 ute=-1.3857143 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12496714 voffcv=0.005 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_3' w0=5e-007 wags=1.9131429e-009 walpha0=6.6315429e-012 wbeta0=8.2628571e-008 wint=1e-008 wk2=-7.1987657e-009 wketa=-9.3497143e-010 wkt1=-5.904e-009 wkt2=1.7142857e-010 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=6.8777143e-009 wr=1 wtvoff=0 wu0=8.1565714e-010 wua=8.016e-018 wub1=3.456e-026 wub=-2.7222857e-026 wuc=-8.7572571e-018 wute=1.7142857e-008 wvoff=2.0674286e-009 wvth0=-1.0069714e-008 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.4 nmos a0=0.10680558 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.35500309 alpha0=2.6500109e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=20.982852 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0036363636 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95938091 k2=0.041255727 k3=0 k3b=0 keta=-0.12490989 kt1=-0.37773746 kt1l=0 kt2=-0.014603854 ku0=0 kvsat=0 kvth0=0 la0=-1.6983636e-009 lags=-1.1780546e-008 lalpha0=-2.8170545e-013 lbeta0=-8.9454546e-008 ldelta=3.1818182e-009 level=54 lint=0 lk1=-9.9985454e-008 lk2=-3.7879164e-008 lketa=3.0254945e-008 lkt1=1.6718727e-008 lkt2=-3.3230727e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=-8.0088e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.0251818e-009 lua=3.9938436e-016 lub1=2.4878e-025 lub=-9.0230909e-026 luc=-3.4349127e-017 lvoff=-9.2114546e-009 lvsat=0.0042909091 lvth0=-4.1979273e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.0504145e-015 pags=-1.3815011e-014 palpha0=-2.4870109e-020 paramchk=1 pbeta0=1.0555636e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.45921829 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=3.5791331e-015 pketa=1.6899316e-015 pkt1=3.5425745e-015 pkt2=1.9005294e-015 ppclm=2.4308858e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.5013818e-016 pua=3.8566691e-024 pub1=-3.8927127e-032 pub=-2.4352626e-031 puc=-7.5187026e-024 pvag=0 pvoff=4.8246982e-015 pvsat=-2.0596364e-009 pvth0=2.0029964e-015 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.033011551 ua1=1.675e-009 ua=-6.3005701e-010 ub1=-3.65896e-018 ub=2.2836418e-018 uc1=-5.6e-011 uc=1.5877203e-010 ute=-1.4342857 vbm=-3 version=4.5 vfbcv=-1 voff=-0.079311948 voffcv=0.005 voffl=0 vsat=71618.182 vth0='nmos_3p3_vth0_4' w0=5e-007 wa0=-3.7514805e-009 wags=3.3067462e-008 walpha0=4.9740218e-014 wbeta0=-3.786053e-007 wint=1e-008 wk2=-1.2782618e-008 wketa=-3.3798633e-009 wkt1=-7.0851491e-009 wkt2=-3.8010589e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.9828414e-008 wr=1 wtvoff=0 wu0=1.2335751e-010 wua=1.8551439e-017 wub1=7.7854254e-026 wub=1.1549411e-025 wuc=-1.9125195e-020 wute=4.0457143e-008 wvoff=-1.7231065e-008 wvsat=0.0097832727 wvth0=-2.1596758e-008 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.5 nmos a0=0.97533082 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.441074 alpha0=6.8164074e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.036008 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0014285714 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.76833212 k2=0.0082103273 k3=0 k3b=0 keta=-0.043888571 kt1=-0.4079911 kt1l=0 kt2=-0.031229592 ku0=0 kvsat=0 kvth0=0 la0=-4.3596098e-007 lags=-5.4816e-008 lalpha0=-2.3649037e-012 lbeta0=-1.1603265e-007 ldelta=4.2857143e-009 level=54 lint=0 lk1=-4.4610612e-009 lk2=-2.1356464e-008 lketa=-1.0255714e-008 lkt1=3.1845551e-008 lkt2=4.9897959e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=4.0921959e-008 lpdiblc2=9.06e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.9403755e-009 lua=6.6367861e-016 lub1=-1.7578531e-025 lub=-3.6042122e-025 luc1=3.1443869e-017 luc=4.0383673e-018 lvoff=1.1378694e-008 lvsat=-0.0041142857 lvth0=-1.7716408e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.4148441e-015 pags=-2.7963977e-014 palpha0=6.6303478e-020 paramchk=1 pbeta0=-2.8990433e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21719837 pdiblc1=0.39 pdiblc2=0.001359 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=5.2640522e-015 pk2=-5.0342094e-015 pkt1=-1.5285865e-014 pkt2=-2.6008163e-015 ppclm=2.4676545e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-3.5579167e-016 pua=2.2512666e-023 pub1=-2.9753339e-032 pub=-2.3455895e-031 puc1=-1.5093057e-023 puc=-9.2762449e-024 pvag=0 pvoff=-6.4985731e-015 pvsat=4.8548571e-009 pvth0=-3.3082384e-015 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.031181163 ua1=1.675e-009 ua=-1.1586455e-009 ub1=-2.8098294e-018 ub=2.8240225e-018 uc1=-1.1888774e-010 uc=8.1997037e-011 ute=-1.4342857 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12049225 voffcv=0.005 voffl=0 vsat=88428.571 vth0='nmos_3p3_vth0_5' w0=5e-007 wa0=1.1790367e-009 wags=6.1365394e-008 walpha0=-1.3260696e-013 wbeta0=4.1231608e-007 wint=1e-008 wk1=-1.0528104e-008 wk2=4.4440669e-009 wkt1=3.0571729e-008 wkt2=5.2016327e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-2.0563788e-008 wr=1 wtvoff=0 wu0=1.3466449e-010 wua=-1.8760555e-017 wub1=5.9506678e-026 wub=9.755951e-026 wuc1=3.0186115e-017 wuc=3.4959595e-018 wute=4.0457143e-008 wvoff=5.4154776e-009 wvsat=-0.0040457143 wvth0=-1.0974289e-008 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.6 nmos a0=1.2333595 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.28370796 alpha0=9.0921047e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.039866 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027272727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79418892 k2=-0.0057236965 k3=0 k3b=0 keta=-0.021025909 kt1=-0.33923366 kt1l=0 kt2=-0.021803571 ku0=0 kvsat=0 kvth0=0 la0=-7.4559545e-007 lags=1.3402325e-007 lalpha0=-1.0329047e-010 lbeta0=-3.7206623e-006 ldelta=2.7272727e-009 level=54 lint=0 lk1=-3.5489221e-008 lk2=-4.6356351e-009 lketa=-3.7690909e-008 lkt1=-5.0663377e-008 lkt2=-6.3214286e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lpclm=2.9060649e-008 lpdiblc2=1.7686364e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=-1.4308442e-009 lua=2.1903156e-016 lub1=7.0824935e-025 lub=-6.4298182e-025 luc1=-5.0024338e-017 luc=-1.4633922e-017 lute=3.448052e-007 lvoff=1.3159091e-008 lvth0=1.325026e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=6.3697932e-014 palpha0=-1.0548281e-019 paramchk=1 pbeta0=-2.9791169e-014 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.22708279 pdiblc1=0.39 pdiblc2=0.00064013636 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-8.3746286e-015 pk2=2.7051485e-015 pkt1=2.4318421e-014 pkt2=3.0342857e-015 ppclm=1.9242888e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=1.3295688e-015 pua=8.5070338e-024 pub1=-5.7827969e-031 pub=8.4187636e-032 puc1=2.4011682e-023 puc=5.071119e-024 pute=-1.6550649e-013 pvag=0 pvth0=-1.1596488e-014 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.036490513 ua1=1.675e-009 ua=-7.881063e-010 ub1=-3.5465249e-018 ub=3.0594896e-018 uc1=-5.0997566e-011 uc=9.7557278e-011 ute=-1.7216234 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12197591 voffcv=0.005 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_6' w0=5e-007 wags=-1.501953e-008 walpha0=1.0548281e-014 wbeta0=1.9555512e-007 wint=1e-008 wk1=8.3746286e-010 wk2=-2.005398e-009 wkt1=-2.4318421e-009 wkt2=5.0571429e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.603574e-008 wr=1 wtvoff=0 wu0=-1.2698026e-009 wua=-7.0891948e-018 wub1=5.1661197e-025 wub=-1.6806265e-025 wuc1=-2.4011682e-018 wuc=-8.460177e-018 wute=1.7837922e-007 wvth0=-4.067414e-009 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.7 nmos a0=1.1588 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29711029 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=23.6678 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79064 k2=-0.00618726 k3=0 k3b=0 keta=-0.024795 kt1=-0.3443 kt1l=0 kt2=-0.022435714 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.22998886 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.036347429 ua1=1.675e-009 ua=-7.6620314e-010 ub1=-3.4757e-018 ub=2.9951914e-018 uc1=-5.6e-011 uc=9.6093886e-011 ute=-1.6871429 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.005 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_7' w0=5e-007 wags=-8.6497371e-009 wbeta0=1.92576e-007 wint=1e-008 wk2=-1.7348832e-009 wkt2=8.0914286e-010 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-1.4111451e-008 wr=1 wtvoff=0 wu0=-1.1368457e-009 wua=-6.2384914e-018 wub1=4.58784e-025 wub=-1.5964389e-025 wuc=-7.9530651e-018 wute=1.6182857e-007 wvth0=-5.2270629e-009 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.8 nmos a0=0.10362636 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.2705431 alpha0=2.5953123e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.140586 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0036363636 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95060511 k2=0.013945175 k3=0 k3b=0 keta=-0.12424077 kt1=-0.28115299 kt1l=0 kt2=-0.025449687 ku0=0 kvsat=0 kvth0=0 la0=-8.0818182e-010 lags=3.2753448e-008 lalpha0=-2.5435614e-013 ldelta=3.1818182e-009 level=54 lint=0 lk1=-9.5597554e-008 lk2=-3.0232209e-008 lketa=2.9920384e-008 lkt1=-1.0099496e-008 lkt2=9.6575269e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.2990496e-006 lpclm=-9.798626e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.7050207e-010 lua=2.5458994e-016 lub1=4.827456e-025 lub=-3.3240512e-025 luc1=4.973267e-017 luc=-6.8059408e-017 lvoff=6.8691116e-010 lvoffcv=-1.118626e-007 lvsat=-0.00034132231 lvth0=-5.5747725e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.59809917 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pags=-6.6365124e-014 palpha0=-5.7142305e-020 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.20476889 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=-5.177723e-015 pk2=-5.4442735e-015 pketa=2.0847148e-015 pkt1=3.5188078e-014 pkt2=-3.1602845e-015 pnoff=-1.5328785e-012 ppclm=-5.8632603e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=4.1983839e-015 pua=1.7471409e-022 pub1=-3.1500653e-031 pub=4.2239319e-032 puc1=-5.8684551e-023 puc=3.2259428e-023 pvag=0 pvoff=-6.8553733e-015 pvoffcv=1.3199787e-013 pvsat=3.4063967e-009 pvth0=1.824977e-014 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.046898182 ua1=1.675e-009 ua=-6.6207759e-010 ub1=-5.3788142e-018 ub=3.7962141e-018 uc1=-2.2938539e-010 uc=2.9436835e-010 ute=-1.5701136 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12424632 voffcv=0.22872521 voffl=0 vsat=85682.645 vth0='nmos_3p3_vth0_8' w0=5e-007 wags=1.3273025e-007 walpha0=1.1428461e-013 wbeta0=-5.6473191e-007 wint=1e-008 wk1=1.0355446e-008 wk2=1.9443834e-008 wketa=-4.1694295e-009 wkt1=-1.2105482e-007 wkt2=8.9970236e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=3.065757e-006 wpclm=2.8042187e-007 wr=1 wtvoff=0 wu0=-1.6262868e-008 wua=5.6335718e-017 wub1=2.1072821e-024 wub=-1.6693412e-024 wuc1=2.0459475e-016 wuc=-1.6002278e-016 wute=2.0073409e-007 wvoff=3.5791497e-008 wvoffcv=-2.6399574e-007 wvsat=-0.0068127934 wvth0=-5.7737207e-008 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.9 nmos a0=0.57970277 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.63340774 alpha0=6.7040286e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.043581 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0014285714 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.017155231 k3=0 k3b=0 keta=-0.043888571 kt1=-0.30297354 kt1l=0 kt2=-0.021799026 ku0=0 kvsat=0 kvth0=0 la0=-2.3884638e-007 lags=-1.4867887e-007 lalpha0=-2.3087143e-012 lbeta0=4.8502597e-008 ldelta=4.2857143e-009 level=54 lint=0 lk2=-3.1837237e-008 lketa=-1.0255714e-008 lkt1=8.1077922e-010 lkt2=-8.5957792e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=6.8726318e-008 lpdiblc2=9.06e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.387089e-009 lua=3.880134e-016 lub1=-6.899552e-025 lub=-1.7056325e-025 luc1=7.5986727e-018 luc=5.1261039e-019 lvoff=-1.0167857e-008 lvth0=-9.953513e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.3401007e-013 pags=8.279421e-014 paramchk=1 pbeta0=-4.8405592e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.047719 pdiblc1=0.39 pdiblc2=0.001359 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk2=7.3331031e-015 pkt1=2.1335166e-014 pkt2=4.3014448e-015 ppclm=-8.1325983e-015 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=2.9708645e-016 pua=3.4779762e-022 pub1=5.7696713e-031 pub=-4.5859137e-031 puc1=1.3044275e-023 puc=-5.1158517e-024 pvag=0 pvoff=1.8926357e-014 pvth0=-1.2468455e-014 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.038465008 ua1=1.675e-009 ua=-9.289245e-010 ub1=-3.0334126e-018 ub=3.4725304e-018 uc1=-1.4511739e-010 uc=1.5722431e-010 ute=-1.5701136 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10253679 voffcv=0.005 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_9' w0=5e-007 wa0=4.6802014e-007 wags=-1.6558842e-007 wbeta0=4.0337993e-007 wint=1e-008 wk2=-6.1109193e-009 wkt1=-9.3348999e-008 wkt2=-5.9264351e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.7942187e-007 wr=1 wtvoff=0 wu0=-8.4602728e-009 wua=-2.8983135e-016 wub1=3.2333483e-025 wub=-6.6767982e-025 wuc1=6.1137104e-017 wuc=-8.5272224e-017 wute=2.0073409e-007 wvoff=-1.5771964e-008 wvth0=3.6992425e-009 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.10 nmos a0=1.175342 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26729169 alpha0=9.0929986e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.512311 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027272727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79747612 k2=-0.0074231864 k3=0 k3b=0 keta=-0.021025909 kt1=-0.31506405 kt1l=0 kt2=-0.016812862 ku0=0 kvsat=0 kvth0=0 la0=-9.536135e-007 lags=2.9066039e-007 lalpha0=-1.0337986e-010 lbeta0=-4.1139731e-006 ldelta=2.7272727e-009 level=54 lint=0 lk1=-4.5679339e-008 lk2=-2.3431364e-009 lketa=-3.7690909e-008 lkt1=1.5319401e-008 lkt2=-6.8429752e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.5464876e-007 lpclm=-1.5414418e-007 lpdiblc2=1.7686364e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.9522345e-009 lua1=2.5980992e-017 lua=2.4617513e-016 lub1=-1.7520434e-024 lub=1.6897655e-025 luc1=-1.1288886e-016 luc=6.3987831e-017 lute=-2.7427686e-008 lvoff=1.3159091e-008 lvoffcv=8.5056818e-008 lvth0=7.3817355e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.128874 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=2.454613e-013 pags=-1.211339e-013 paramchk=1 pbeta0=4.3431558e-013 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23344442 pdiblc1=0.39 pdiblc2=0.00064013636 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pk1=3.6497107e-015 pkt1=-5.3541257e-014 pkt2=3.6497107e-015 pnoff=1.8248554e-013 ppclm=2.3542459e-013 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pu0=-2.662464e-015 pua1=-3.065757e-023 pua=-2.3522386e-023 pub1=2.3248657e-030 pub=-8.7392324e-031 puc1=9.8191818e-023 puc=-8.7702549e-023 pute=2.7372831e-013 pvag=0 pvoffcv=-1.0036705e-013 pvth0=-4.6716298e-015 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040494054 ua1=1.6533492e-009 ua=-8.1072595e-010 ub1=-2.1483391e-018 ub=3.1895805e-018 uc1=-4.4711114e-011 uc=1.0432829e-010 ute=-1.5472572 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12197591 voffcv=-0.065880682 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_10' w0=5e-007 wa0=6.8460666e-008 wags=4.3516718e-009 wbeta0=-3.6192965e-007 wint=1e-008 wk1=-3.0414256e-009 wkt1=-3.095198e-008 wkt2=-5.3833233e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.5207128e-007 wpclm=-2.3542459e-008 wr=1 wtvoff=0 wu0=-5.9939808e-009 wua1=2.5547975e-017 wua=1.9601988e-017 wub1=-1.1332474e-024 wub=-3.2156993e-025 wuc1=-9.8191818e-018 wuc=-1.6449976e-017 wute=-2.7372831e-008 wvoffcv=8.3639205e-008 wvth0=-2.7981116e-009 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.11 nmos a0=1.0799807 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29635773 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.100914 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79290818 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31353211 kt1l=0 kt2=-0.017497159 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1134091 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040689277 ua1=1.6559473e-009 ua=-7.8610843e-010 ub1=-2.3235434e-018 ub=3.2064782e-018 uc1=-5.6e-011 uc=1.1072708e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.057375 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_11' w0=5e-007 wa0=9.3006796e-008 wags=-7.7617182e-009 wbeta0=-3.1849809e-007 wint=1e-008 wk1=-2.6764545e-009 wkt1=-3.6306106e-008 wkt2=-5.0183523e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wnoff=-1.3382273e-007 wr=1 wtvoff=0 wu0=-6.2602272e-009 wua1=2.2482218e-017 wua=1.7249749e-017 wub1=-9.0076078e-025 wub=-4.0896225e-025 wuc=-2.5220231e-017 wvoffcv=7.36025e-008 wvth0=-3.2652745e-009 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.12 nmos a0=0.13211844 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.46155061 alpha0=2.6067636e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=2.3e-010 cgidl=0.5 cgsl=1e-010 cgso=2.3e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0036363636 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.95164273 k2=0.015893454 k3=0 k3b=0 keta=-0.12105603 kt1=-0.29328273 kt1l=0 kt2=-0.024548182 ku0=0 kvsat=0 kvth0=0 la0=-1.5054221e-008 lags=-6.2750307e-008 lalpha0=-2.6008182e-013 ldelta=3.1818182e-009 level=54 lint=0 lk1=-9.6116364e-008 lk2=-3.0777727e-008 lketa=2.8328017e-008 lkt1=-6.5736364e-009 lkt2=6.4909091e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lnoff=1.1454545e-006 lpclm=-1.5673636e-008 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=5.9118182e-010 lua=2.7209636e-016 lub1=4.5118182e-025 lub=-3.2817273e-025 luc1=4.3852454e-017 luc=-6.4827e-017 lvoffcv=-9.8636364e-008 lvth0=-5.3919091e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=-0.29090909 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=1.4217547e-013 pags=8.8676235e-013 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23286727 pdiblc1=0.39 pdiblc2=0.003171 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 pketa=1.7976533e-014 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.045268636 ua1=1.675e-009 ua=-6.5643273e-010 ub1=-5.1676636e-018 ub=3.6289455e-018 uc1=-2.0888491e-010 uc=2.78334e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=0.20227273 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_12' w0=5e-007 wa0=-2.8435094e-007 wags=-1.7735247e-006 wint=1e-008 wketa=-3.5953066e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.13 nmos a0=0.62659857 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.61681571 alpha0=6.7040286e-006 alpha1=0 at=23000 b0=0 b1=0 beta0=21.084 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0014285714 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.75941 k2=0.016542914 k3=0 k3b=0 keta=-0.043888571 kt1=-0.31232714 kt1l=0 kt2=-0.022392857 ku0=0 kvsat=0 kvth0=0 la0=-2.6229429e-007 lags=-1.4038286e-007 lalpha0=-2.3087143e-012 ldelta=4.2857143e-009 level=54 lint=0 lk2=-3.1102457e-008 lketa=-1.0255714e-008 lkt1=2.9485714e-009 lkt2=-4.2857143e-010 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=6.7911429e-008 lpdiblc2=9.06e-010 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=4.4168571e-009 lua=4.2286286e-016 lub1=-6.3214286e-025 lub=-2.1651429e-025 luc1=8.9057143e-018 lvoff=-8.2714286e-009 lvth0=-1.1202857e-008 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.065697143 pdiblc1=0.39 pdiblc2=0.001359 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.037617286 ua1=1.675e-009 ua=-9.5796571e-010 ub1=-3.0010143e-018 ub=3.4056286e-018 uc1=-1.3899143e-010 uc=1.4868e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.10411714 voffcv=0.005 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_13' w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.14 nmos a0=1.1822018 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.26772773 alpha0=9.0929986e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.476046 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=1e-010 cgidl=0.5 cgsl=1e-010 cgso=1e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.0027272727 diomod=1 dlc=0 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79717136 k2=-0.0074231864 k3=0 k3b=0 keta=-0.021025909 kt1=-0.31816545 kt1l=0 kt2=-0.017352273 ku0=0 kvsat=0 kvth0=0 la0=-9.2901818e-007 lags=2.7852273e-007 lalpha0=-1.0337986e-010 lbeta0=-4.0704545e-006 ldelta=2.7272727e-009 level=54 lint=0 lk1=-4.5313636e-008 lk2=-2.3431364e-009 lketa=-3.7690909e-008 lkt1=9.9545454e-009 lkt2=-6.4772727e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=-1.3636364e-007 lpclm=-1.3055455e-007 lpdiblc2=1.7686364e-009 lpe0=1.1e-007 lpeb=0 ltvoff=0 lu0=1.6854546e-009 lua1=2.2909091e-017 lua=2.4381818e-016 lub1=-1.5190909e-024 lub=8.1409091e-026 luc1=-1.0305e-016 luc=5.52e-017 lvoff=1.3159091e-008 lvoffcv=7.5e-008 lvth0=6.9136364e-009 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1136364 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.23108545 pdiblc1=0.39 pdiblc2=0.00064013636 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.039893455 ua1=1.6559091e-009 ua=-8.0876182e-010 ub1=-2.2618909e-018 ub=3.1573591e-018 uc1=-4.5695e-011 uc=1.0268e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12197591 voffcv=-0.0575 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_14' w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.model nmos_3p3.15 nmos a0=1.0893 a1=0 a2=1 acde=0.6 acnqsmod=0 agidl=1.3268e-010 ags=0.29558 alpha0=8.0592e-005 alpha1=0 at=23000 b0=0 b1=0 beta0=24.069 bgidl=1.8961e+009 binunit=2 capmod=2 cdsc=0 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=1e-010 cgdo=2.3e-010 cgidl=0.5 cgsl=1e-010 cgso=2.3e-010 cit=0 cjs=0.00096797 cjswgs=5.9903e-010 cjsws=1.5663e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.003 diomod=1 dlc=3e-008 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.5 dvt0=0 dvt0w=0 dvt1=0.53 dvt1w=0 dvt2=0 dvt2w=0 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=0.95 egidl=0.8 em=4.1e+007 epsrox=3.9 eta0=0.75 etab=-0.32 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=2.2959e-007 jswgs=0 jsws=2.1207e-013 k1=0.79264 k2=-0.0076575 k3=0 k3b=0 keta=-0.024795 kt1=-0.31717 kt1l=0 kt2=-0.018 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=1.1e-007 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.25 mjs=0.32071 mjswgs=0.32059 mjsws=0.1 mobmod=0 moin=15 ndep=3e+017 nfactor=1 ngate=6e+019 njs=1.01 noff=2.1 noia='nmos_3p3_noia' noib='nmos_3p3_noib' noic='nmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.70172 pbswgs=0.74743 pbsws=0.8062 pclm=0.21803 pdiblc1=0.39 pdiblc2=0.000817 pdiblcb=0.2 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.07 prt=0 prwb=0 prwg=0 pscbe1=6.6469e+008 pscbe2=1.638e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='nmos_3p3_rdsw' rdswmin=50 rdwmin=0 rgatemod=0 rsh=7 rswmin=0 saref=4.4e-007 sbref=4.4e-007 tcj=0.0009438 tcjsw=0.00060474 tcjswg=0.001 tnoimod=0 tnom=25 toxe='nmos_3p3_tox' toxm=8e-009 toxp='nmos_3p3_tox' toxref=8e-009 tpb=0.0018129 tpbsw=5e-005 tpbswg=0.0016872 trnqsmod=0 tvoff=0.001 u0=0.040062 ua1=1.6582e-009 ua=-7.8438e-010 ub1=-2.4138e-018 ub=3.1655e-018 uc1=-5.6e-011 uc=1.082e-010 ute=-1.55 vbm=-3 version=4.5 vfbcv=-1 voff=-0.12066 voffcv=-0.05 voffl=0 vsat=85000 vth0='nmos_3p3_vth0_15' w0=5e-007 wint=1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wr=1 wtvoff=0 ww=0 wwl=0 wwn=1 xj='nmos_3p3_xj' xl='nmos_3p3_xl' xpart=0 xtis=3 xw='nmos_3p3_xw'
.subckt nplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 r_rsh0='rsh_nplus_u_m' r_dw=-5e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.36e-3 r_tc2=6.5e-7 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model np_junction d cj=0.00096797 level=2
d1 3 1 np_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends nplus_u_m1
.endl nmos_3p3_stat

.lib pmos_3p3_stat
.subckt pmos_3p3_sab d g s b w=10u l=0.28u par=1 s_sab=0.48u d_sab=1.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.00666
.param par_k=0.002833
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b pplus_u_m1 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b pplus_u_m1 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b pmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='sa' sb='sb' sd='sd' delvto='mis_vth*sw_stat_mismatch'
.ends
.model pmos_3p3.0 pmos a0=1.0272635 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19081247 alpha0=1.1485698e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=39.773597 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.86959286 k2=0.029351195 k3=0 k3b=0 keta=-0.066404636 kt1=-0.28373805 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.0434818e-007 lags=1.0492091e-007 lalpha0=-3.0054064e-012 lbeta0=-3.6237273e-006 level=54 lint=0 lk1=4.91e-009 lk2=-2.4890454e-008 lketa=8.2658182e-009 lkt1=-1.5974545e-008 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=7.0823636e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.4492727e-009 lua1=1.7181818e-016 lua=1.0386891e-015 lub1=-6.7359091e-025 lub=-1.4361909e-025 luc1=5.8570909e-017 luc=8.4861818e-018 lvoff=-1.6014546e-009 lvth0=-7.6827273e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-2.7370909e-015 pags=-1.2080073e-014 palpha0=6.39288e-020 paramchk=1 pbeta0=1.1827636e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.35627558 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-2.0974909e-014 pk2=3.4158327e-015 pketa=3.6614618e-015 pkt1=1.9400727e-015 ppclm=6.5406545e-015 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-5.2642909e-016 pua1=-8.9345454e-023 pua=-1.9180342e-022 pub1=1.4950473e-031 pub=1.3557818e-033 puc1=-1.4057018e-023 puc=-4.4743636e-024 pvag=0 pvoff=8.3275636e-016 pvth0=2.3570182e-015 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0077071688 ua1=1.1563636e-009 ua=-2.4381818e-012 ub1=-2.100161e-018 ub=6.7035533e-019 uc1=-2.5418182e-010 uc=8.6801065e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094658091 voffcv=-0.16 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_0' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.1112467e-008 wags=-2.3219283e-008 walpha0=-1.0325417e-013 wbeta0=2.1005299e-007 wint=-1e-008 wk1=6.7137132e-008 wk2=-2.1522854e-008 wketa=-7.3229236e-009 wkt1=-1.1172031e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=2.9266005e-008 wtvoff=0 wu0=6.0892675e-010 wua1=1.7869091e-016 wua=3.3100364e-018 wub1=-1.4002317e-025 wub=-4.8420779e-027 wuc1=4.0843636e-017 wuc=-1.3364176e-017 wvoff=-1.6655127e-009 wvth0=4.2938493e-009 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.1 pmos a0=1.1510659 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19022326 alpha0=7.5504633e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=42.422959 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.011648 k2=-0.018784 k3=0 k3b=0 keta=-0.0050909592 kt1=-0.30703735 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.6624939e-007 lags=1.0521551e-007 lalpha0=-3.5014873e-011 lbeta0=-4.9484082e-006 level=54 lint=0 lk1=-6.6117551e-008 lk2=-8.2285714e-010 lketa=-2.239102e-008 lkt1=-4.324898e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=1.2067592e-007 lpdiblc2=2.4533143e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.1587837e-009 lua=8.5199265e-016 lub1=-6.0410204e-025 lub=-3.5234082e-025 luc1=-3.0738122e-017 luc=5.8519641e-017 lvoff=1.2890571e-008 lvth0=8.0902041e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.6645518e-014 pags=-3.0616751e-014 palpha0=-2.3899709e-018 paramchk=1 pbeta0=8.5195102e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.25657102 pdiblc1=0.1484 pdiblc2=0.00024628714 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=2.1589126e-014 pk2=-6.084e-015 pketa=1.1021878e-015 pkt1=-1.6167967e-014 ppclm=-2.1505078e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-9.8910367e-017 pua=-1.6858315e-022 pub1=9.6045061e-032 pub=9.5112882e-032 puc1=3.2542237e-024 puc=-7.4630909e-024 pvag=0 pvth0=1.5205225e-015 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010288147 ua1=1.5e-009 ua=3.7095469e-010 ub1=-2.2391388e-018 ub=1.0877988e-018 uc1=-7.5563755e-011 uc=-1.3265853e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12364214 voffcv=-0.16 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_1' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=3.8929322e-008 wags=1.3854074e-008 walpha0=4.8045453e-012 wbeta0=2.7621551e-007 wint=-1e-008 wk1=-1.7990939e-008 wk2=-2.5231886e-009 wketa=-2.2043755e-009 wkt1=2.5044049e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=8.5357469e-008 wtvoff=0 wu0=-2.4611069e-010 wua=-4.3130498e-017 wub1=-3.3103837e-026 wub=-1.9235628e-025 wuc1=6.2211526e-018 wuc=-7.386721e-018 wvth0=5.9668408e-009 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.2 pmos a0=1.2626103 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.15731682 alpha0=0.0020588939 alpha1=0 at=12000 b0=0 b1=0 beta0=44.45026 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95493474 k2=-0.010993416 k3=0 k3b=0 keta=-0.00016272403 kt1=-0.26850506 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-4.001026e-007 lags=1.4470325e-007 lalpha0=-2.415082e-009 lbeta0=-7.3811688e-006 level=54 lint=0 lk1=1.9383117e-009 lk2=-1.0171558e-008 lketa=-2.8304903e-008 lkt1=-5.0563636e-008 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4545454e-007 lpclm=4.2841558e-008 lpdiblc2=4.4675455e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=3.0025909e-009 lua=8.1926494e-016 lub1=3.3323377e-025 lub=-6.9161688e-026 luc1=-7.8734805e-017 luc=9.5515247e-017 lvoff=-1.8220325e-008 lvoffcv=-2.1818182e-007 lvth0=-9.5551948e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9454546 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=3.4170078e-014 pags=-1.4866597e-014 palpha0=-2.3332535e-017 paramchk=1 pbeta0=-6.7464935e-014 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32143299 pdiblc1=0.1484 pdiblc2=7.8434545e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk1=-3.6710649e-014 pk2=8.9552104e-015 pketa=2.6125948e-015 pkt1=2.6293091e-014 ppclm=7.4952935e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-6.5690182e-016 pua=-1.5714468e-022 pub1=-1.7328156e-031 pub=-4.1208312e-033 puc1=2.5455553e-023 puc=-1.8553586e-023 pvag=0 pvoff=-1.1894494e-015 pvth0=4.2667013e-015 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0087516409 ua1=1.5e-009 ua=3.9822779e-010 ub1=-3.0202519e-018 ub=8.5181617e-019 uc1=-3.5566519e-011 uc=-4.4095525e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097716396 voffcv=0.021818182 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_2' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-3.4170078e-009 wags=7.2894545e-010 walpha0=2.2256682e-011 wbeta0=4.0343221e-007 wint=-1e-008 wk1=3.0592208e-008 wk2=-1.5055864e-008 wketa=-3.463048e-009 wkt1=-1.0340166e-008 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=4.9757922e-009 wtvoff=0 wu0=2.1888218e-010 wua=-5.2662561e-017 wub1=1.9133501e-025 wub=-1.0966152e-025 wuc1=-1.2279955e-017 wuc=1.8553586e-018 wvoff=9.9120779e-010 wvth0=3.6783584e-009 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.3 pmos a0=1.2226 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17178714 alpha0=0.0018173857 alpha1=0 at=12000 b0=0 b1=0 beta0=43.712143 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.95512857 k2=-0.012010571 k3=0 k3b=0 keta=-0.0029932143 kt1=-0.27356143 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32571714 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0090519 ua1=1.5e-009 ua=4.8015429e-010 ub1=-2.9869286e-018 ub=8.449e-019 uc1=-4.344e-011 uc=-3.4544e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.099538429 voffcv=0 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_3' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-7.5771429e-010 walpha0=1.9923429e-011 wbeta0=3.9668571e-007 wint=-1e-008 wk1=2.6921143e-008 wk2=-1.4160343e-008 wketa=-3.2017886e-009 wkt1=-7.7108571e-009 wl=0 wln=1 wmax=5e-007 wmin=2.2e-007 wpclm=1.2471086e-008 wtvoff=0 wu0=1.53192e-010 wua=-6.8377029e-017 wub1=1.7400686e-025 wub=-1.100736e-025 wuc1=-9.7344e-018 wvoff=8.7226286e-010 wvth0=4.1050286e-009 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.4 pmos a0=0.66833429 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20459958 alpha0=1.2079775e-005 alpha1=0 at=12000 b0=0 b1=0 beta0=38.238696 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99870273 k2=0.014249873 k3=0 k3b=0 keta=-0.10490303 kt1=-0.33225761 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-1.03128e-007 lags=6.9689636e-008 lalpha0=-3.0255502e-012 lbeta0=-2.7152909e-006 level=54 lint=0 lk1=-3.5426364e-008 lk2=-2.0467636e-008 lketa=2.2143527e-008 lkt1=5.3309091e-010 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=2.7248545e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.8372909e-009 lua1=-2.562e-016 lua=7.4813818e-016 lub1=-2.9730909e-026 lub=-3.0903909e-025 luc1=-3.4608e-017 luc=1.2453182e-017 lvth0=-2.1407273e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-5.5371585e-014 pags=6.2401891e-015 palpha0=7.4403585e-020 paramchk=1 pbeta0=-3.5411055e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3781492 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=1.1159673e-015 pketa=-3.5549469e-015 pkt1=-6.6438982e-015 ppclm=2.9199702e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-2.0819854e-016 pua1=1.33224e-022 pua=-4.0716945e-023 pub1=-1.8530247e-031 pub=8.7374182e-032 puc1=3.4396015e-023 puc=-6.5372036e-024 pvag=0 pvth0=-5.2482182e-016 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0091928468 ua1=2.0124e-009 ua=-8.0522078e-011 ub1=-2.8876353e-018 ub=1.748897e-018 uc1=6.432e-012 uc=8.6704408e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_4' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.9775566e-007 wags=-3.0388584e-008 walpha0=-4.121738e-013 wbeta0=1.0082017e-006 wint=-1e-008 wk2=-1.3670166e-008 wketa=1.2696239e-008 wkt1=1.4058139e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.7891728e-008 wtvoff=0 wu0=-1.6362577e-010 wua1=-2.66448e-016 wua=4.3913662e-017 wub1=2.6946346e-025 wub=-5.6568377e-025 wuc1=-9.4675549e-017 wuc=-1.3313914e-017 wvth0=1.4897689e-008 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.5 pmos a0=1.3454526 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.19226653 alpha0=0.000123026 alpha1=0 at=12000 b0=0 b1=0 beta0=43.366204 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.97705 k2=-0.026847376 k3=0 k3b=0 keta=-0.0016565918 kt1=-0.28366163 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-4.4168718e-007 lags=7.5856163e-008 lalpha0=-5.8498663e-011 lbeta0=-5.2790449e-006 level=54 lint=0 lk1=-2.46e-008 lk2=8.0987755e-011 lketa=-2.947969e-008 lkt1=-2.3764898e-008 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=-5.9909388e-008 lpdiblc2=2.4533143e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.5601469e-009 lua=5.7398498e-016 lub1=9.5240816e-026 lub=-7.120898e-026 luc1=1.8185143e-017 luc=5.1804544e-017 lvoff=1.2890571e-008 lvth0=-3.242449e-010 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.4582136e-014 pags=-1.5349891e-014 palpha0=9.8215995e-018 paramchk=1 pbeta0=2.571262e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.55246506 pdiblc1=0.1484 pdiblc2=0.00024628714 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-6.5539994e-015 pketa=4.7882958e-015 pkt1=-6.0591673e-015 ppclm=7.2399282e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-3.0761926e-016 pua=-2.4019161e-023 pub1=-2.6761322e-031 pub=-5.1075673e-032 puc1=-2.2185874e-023 puc=-3.9712404e-024 pvag=0 pvth0=5.8960359e-015 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097471347 ua1=1.5e-009 ua=2.6778433e-010 ub1=-3.1375788e-018 ub=1.2732368e-018 uc1=-9.9154286e-011 uc=8.0016841e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.12364214 voffcv=-0.16 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_5' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-6.215178e-008 wags=1.2791576e-008 walpha0=-1.9906566e-011 wbeta0=-2.1427184e-007 wint=-1e-008 wk2=1.6697667e-009 wketa=-3.9902465e-009 wkt1=1.2888678e-008 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=-6.8507432e-008 wtvoff=0 wu0=3.5215673e-011 wua=1.0518093e-017 wub1=4.3408496e-025 wub=-2.8878406e-025 wuc1=1.8488229e-017 wuc=-1.844584e-017 wvth0=2.0559739e-009 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.6 pmos a0=1.1189871 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16561084 alpha0=0.002173683 alpha1=0 at=12000 b0=0 b1=0 beta0=44.354662 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0137659 k2=-0.027452061 k3=0 k3b=0 keta=-0.0068224318 kt1=-0.33774851 kt1l=0 kt2=-0.016947818 ku0=0 kvsat=0 kvth0=0 la0=-1.6992857e-007 lags=1.0784299e-007 lalpha0=-2.519287e-009 lbeta0=-6.4651948e-006 level=54 lint=0 lk1=-6.8659091e-008 lk2=8.0661039e-010 lketa=-2.3280682e-008 lkt1=4.1139351e-008 lkt2=4.6581818e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4545454e-007 lpclm=2.0841896e-007 lpdiblc2=4.4675455e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.5779454e-009 lua=4.1154156e-016 lub1=-5.5351558e-025 lub=5.7264156e-026 luc1=-4.9745455e-017 luc=6.0010667e-017 lvoff=-2.0507727e-008 lvoffcv=-2.1818182e-007 lvth0=-1.3737662e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9454546 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-8.5520416e-014 pags=4.3007377e-015 palpha0=3.0854085e-017 paramchk=1 pbeta0=-5.4377143e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3288581 pdiblc1=0.1484 pdiblc2=7.8434545e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=3.2465626e-015 pkt1=-2.1392462e-014 pkt2=-2.4222546e-015 ppclm=-1.1147314e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=8.3913818e-017 pua=5.487148e-023 pub1=2.878281e-031 pub=-6.986227e-032 puc1=1.0381091e-023 puc=-9.1205299e-026 pvag=0 pvth0=1.2358442e-017 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0097323026 ua1=1.5e-009 ua=4.0315384e-010 ub1=-2.5969484e-018 ub=1.1661759e-018 uc1=-4.2545455e-011 uc=1.1632475e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.095810227 voffcv=0.021818182 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_6' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=7.1267013e-008 wags=-3.583948e-009 walpha0=-3.7433637e-011 wbeta0=4.5314286e-007 wint=-1e-008 wk2=-6.4973683e-009 wkt1=2.5666423e-008 wkt2=2.0185455e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wpclm=1.1147314e-009 wtvoff=0 wu0=-2.910619e-010 wua=-5.5224108e-017 wub1=-2.878281e-026 wub=-2.7312856e-025 wuc1=-8.6509091e-018 wuc=-2.1679203e-017 wvth0=6.9590384e-009 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.7 pmos a0=1.1019943 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17639514 alpha0=0.0019217543 alpha1=0 at=12000 b0=0 b1=0 beta0=43.708143 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.0273714 k3=0 k3b=0 keta=-0.0091505 kt1=-0.33363457 kt1l=0 kt2=-0.016482 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.0098900971 ua1=1.5e-009 ua=4.44308e-010 ub1=-2.6523e-018 ub=1.1719023e-018 uc1=-4.752e-011 uc=7.1643143e-012 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_7' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=6.2714971e-008 wags=-3.1538743e-009 walpha0=-3.4348229e-011 wbeta0=3.9876571e-007 wint=-1e-008 wk2=-6.172712e-009 wkt1=2.3527177e-008 wkt2=1.77632e-009 wl=0 wln=1 wmax=1.2e-006 wmin=5e-007 wtvoff=0 wu0=-2.8267051e-010 wua=-4.973696e-017 wub=-2.8011479e-025 wuc1=-7.6128e-018 wuc=-2.1688323e-017 wvth0=6.9602743e-009 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.8 pmos a0=0.8879706 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.3341873 alpha0=9.723125e-006 alpha1=0 at=12000 b0=0 b1=0 beta0=37.805966 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99870273 k2=-0.00067810868 k3=0 k3b=0 keta=-0.088919542 kt1=-0.29596713 kt1l=0 kt2=-0.020842369 ku0=0 kvsat=0 kvth0=0 la0=-1.4725376e-007 lags=-2.4436508e-009 lalpha0=-2.2830898e-012 lbeta0=-2.3737058e-006 level=54 lint=0 lk1=-3.5426364e-008 lk2=-1.7691446e-008 lketa=1.7668152e-008 lkt1=-8.3979897e-009 lkt2=2.1773833e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=5.0559583e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.7890915e-009 lua1=-1.5583996e-016 lua=6.3071157e-016 lub1=-1.2857843e-025 lub=3.2915171e-026 luc1=8.8928926e-019 luc=-7.439668e-018 lvth0=-8.7733719e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.5381528e-015 pags=9.42428e-014 palpha0=-8.3139811e-019 paramchk=1 pbeta0=-7.708444e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.32482036 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-2.2709854e-015 pketa=1.9050111e-015 pkt1=4.2520201e-015 pkt2=-2.6564076e-015 ppclm=7.6023645e-016 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.493953e-016 pua1=1.078475e-023 pua=1.0254352e-022 pub1=-6.4708497e-032 pub=-3.2981002e-031 puc1=-8.9106783e-024 puc=1.7732073e-023 pvag=0 pvth0=7.5670046e-015 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011352976 ua1=1.8116799e-009 ua=3.4788822e-010 ub1=-2.5843988e-018 ub=9.2772209e-019 uc1=-8.5778578e-011 uc=1.3375779e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_8' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-7.0200638e-008 wags=-1.884856e-007 walpha0=2.4629388e-012 wbeta0=1.5361323e-006 wint=-1e-008 wk2=4.5419708e-009 wketa=-6.803611e-009 wkt1=-3.0216242e-008 wkt2=9.4871699e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=8.2952909e-008 wtvoff=0 wu0=-2.7989835e-009 wua1=-2.1569499e-017 wua=-4.7874691e-016 wub1=-1.0048507e-025 wub=4.3614967e-025 wuc1=1.7821357e-017 wuc=-7.0719038e-017 wvth0=4.2305517e-009 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.9 pmos a0=1.1782327 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20788505 alpha0=0.00011108151 alpha1=0 at=12000 b0=0 b1=0 beta0=43.187318 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.97705 k2=-0.030551827 k3=0 k3b=0 keta=-0.0066799724 kt1=-0.30269355 kt1l=0 kt2=-0.010621998 ku0=0 kvsat=0 kvth0=0 la0=-2.9238479e-007 lags=6.0707474e-008 lalpha0=-5.296228e-011 lbeta0=-5.0643818e-006 level=54 lint=0 lk1=-2.46e-008 lk2=-2.7545864e-009 lketa=-2.3451633e-008 lkt1=-5.0347792e-009 lkt2=-2.9328019e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.407763e-008 lpdiblc2=2.4533143e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.4020669e-009 lua=6.4174442e-016 lub1=-1.8989494e-025 lub=1.5676208e-026 luc1=-2.4594545e-017 luc=7.3318673e-017 lvoff=-1.787102e-009 lvth0=-7.1445584e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=-1.0756678e-013 pags=3.1315103e-015 palpha0=3.0672131e-018 paramchk=1 pbeta0=-4.7627532e-015 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.37778426 pdiblc1=0.1484 pdiblc2=0.00024628714 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-3.0945989e-015 pketa=-2.5659333e-015 pkt1=-2.8909912e-014 pkt2=3.5780184e-015 ppclm=-3.006488e-014 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=-1.3347616e-015 pua=-1.0668567e-022 pub1=8.0252392e-032 pub=-1.570756e-031 puc1=3.0005345e-023 puc=-3.0218479e-023 pvag=0 pvoff=1.7906761e-014 pvth0=1.4216818e-014 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010127025 ua1=1.5e-009 ua=3.2582253e-010 ub1=-2.4617658e-018 ub=9.6220002e-019 uc1=-3.4810909e-011 uc=-2.7758895e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.094286796 voffcv=-0.16 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_9' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=1.4185662e-007 wags=-6.2630205e-009 walpha0=-5.3342836e-012 wbeta0=3.968961e-009 wint=-1e-008 wk2=6.1891978e-009 wketa=2.1382778e-009 wkt1=3.6107623e-008 wkt2=-2.981682e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=1.4460314e-007 wtvoff=0 wu0=-4.282509e-010 wua=-6.0288518e-017 wub1=-3.9040685e-025 wub=9.0680837e-026 wuc1=-6.0010691e-017 wuc=2.5182066e-017 wvoff=-3.5813523e-008 wvth0=-9.069076e-009 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.10 pmos a0=1.1832393 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16685819 alpha0=0.0021426891 alpha1=0 at=12000 b0=0 b1=0 beta0=44.161948 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0137659 k2=-0.036023042 k3=0 k3b=0 keta=-0.0068224318 kt1=-0.29670927 kt1l=0 kt2=-0.012757219 ku0=0 kvsat=0 kvth0=0 la0=-2.9839274e-007 lags=1.0993971e-007 lalpha0=-2.4908914e-009 lbeta0=-6.233938e-006 level=54 lint=0 lk1=-6.8659091e-008 lk2=3.8108709e-009 lketa=-2.3280682e-008 lkt1=-1.2215919e-008 lkt2=-3.7053719e-010 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4545454e-007 lpclm=6.5657665e-008 lpdiblc2=4.4675455e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.3166262e-009 lua1=1.2483595e-016 lua=2.315961e-016 lub1=4.4029649e-026 luc1=1.3542397e-017 luc=5.9935909e-017 lvoff=2.8431167e-009 lvoffcv=-2.1818182e-007 lvth0=-4.4690083e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9454546 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 pa0=7.1205867e-014 pags=1.7427347e-015 palpha0=-3.7885537e-018 paramchk=1 pbeta0=-8.2590471e-013 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34313423 pdiblc1=0.1484 pdiblc2=7.8434545e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 pk2=-4.1863519e-016 pkt1=4.3700967e-014 pkt2=3.7127826e-015 ppclm=1.6302147e-013 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pu0=4.0272326e-016 pua1=-1.5229986e-022 pua=2.7440495e-022 pub1=-4.4117708e-031 puc1=-6.6830088e-023 pvag=0 pvoff=-2.848803e-014 pvth0=3.7885537e-015 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011031559 ua1=1.39597e-009 ua=6.676128e-010 ub1=-2.656703e-018 ub=9.7526352e-019 uc1=-6.6591694e-011 uc=-1.6606591e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.098145312 voffcv=0.021818182 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_10' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wa0=-7.1205867e-009 wags=-5.1057076e-009 walpha0=3.7885537e-013 wbeta0=6.8825393e-007 wint=-1e-008 wk2=3.9592281e-009 wkt1=-2.4401443e-008 wkt2=-3.0939855e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wpclm=-1.6302147e-008 wtvoff=0 wu0=-1.8761549e-009 wua1=1.2691655e-016 wua=-3.7786403e-016 wub1=4.4117708e-026 wub=-4.0215498e-026 wuc1=2.0685503e-017 wvoff=2.848803e-009 wvth0=-3.7885537e-010 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.11 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17785216 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.538555 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035641955 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29793086 kt1l=0 kt2=-0.012794273 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011163222 ua1=1.4084536e-009 ua=6.9077241e-010 ub1=-2.6523e-018 ub=9.7526352e-019 uc1=-6.5237455e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_11' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wags=-4.9314341e-009 wbeta0=6.0566345e-007 wint=-1e-008 wk2=3.9173646e-009 wkt1=-2.0031346e-008 wkt2=-2.7227073e-009 wl=0 wln=1 wmax=1e-005 wmin=1.2e-006 wtvoff=0 wu0=-1.8358826e-009 wua1=1.1168656e-016 wua=-3.5042354e-016 wub=-4.0215498e-026 wuc1=1.4002494e-017 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.12 pmos a0=0.88096455 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.31537636 alpha0=9.9689273e-006 alpha1=0 at=12000 b0=0 b1=0 beta0=37.959273 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.99870273 k2=-0.00022481818 k3=0 k3b=0 keta=-0.089598545 kt1=-0.29898273 kt1l=0 kt2=-0.019895546 ku0=0 kvsat=0 kvth0=0 la0=-1.4740727e-007 lags=6.9618182e-009 lalpha0=-2.3660636e-012 lbeta0=-2.4506364e-006 level=54 lint=0 lk1=-3.5426364e-008 lk2=-1.7918091e-008 lketa=1.7858273e-008 lkt1=-7.9736364e-009 lkt2=1.9122727e-009 ll=0 lln=1 lmax=5e-007 lmin=2.8e-007 lpclm=5.0635454e-008 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.7741818e-009 lua1=-1.5476364e-016 lua=6.4094546e-016 lub1=-1.3503636e-025 luc=-5.67e-018 lvth0=-8.0181818e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.33309909 pdiblc1=0.1484 pdiblc2=0.00073695 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.011073636 ua1=1.8095273e-009 ua=3.0010909e-010 ub1=-2.5944273e-018 ub=9.7125e-019 uc1=-8.4e-011 uc=1.267e-010 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_12' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.13 pmos a0=1.19239 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.20726 alpha0=0.00011054914 alpha1=0 at=12000 b0=0 b1=0 beta0=43.187714 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=0.97705 k2=-0.029934143 k3=0 k3b=0 keta=-0.0064665714 kt1=-0.29909 kt1l=0 kt2=-0.010919571 ku0=0 kvsat=0 kvth0=0 la0=-3.0312e-007 lags=6.102e-008 lalpha0=-5.2656171e-011 lbeta0=-5.0648571e-006 level=54 lint=0 lk1=-2.46e-008 lk2=-3.0634286e-009 lketa=-2.3707714e-008 lkt1=-7.92e-009 lkt2=-2.5757143e-009 ll=0 lln=1 lmax=1.2e-006 lmin=5e-007 lpclm=2.1077143e-008 lpdiblc2=2.4533143e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=2.2688571e-009 lua=6.3109714e-016 lub1=-1.8188571e-025 luc1=-2.16e-017 luc=7.0302857e-017 lvth0=-5.7257143e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2.4 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.39221571 pdiblc1=0.1484 pdiblc2=0.00024628714 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010084286 ua1=1.5e-009 ua=3.1980571e-010 ub1=-2.5007286e-018 ub=9.7125e-019 uc1=-4.08e-011 uc=-2.5245714e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=-0.16 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_13' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.14 pmos a0=1.1825286 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.16634864 alpha0=0.002142727 alpha1=0 at=12000 b0=0 b1=0 beta0=44.230636 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0137659 k2=-0.035627909 k3=0 k3b=0 keta=-0.0068224318 kt1=-0.29914454 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 la0=-2.9128636e-007 lags=1.1011364e-007 lalpha0=-2.4912696e-009 lbeta0=-6.3163636e-006 level=54 lint=0 lk1=-6.8659091e-008 lk2=3.7690909e-009 lketa=-2.3280682e-008 lkt1=-7.8545455e-009 ll=0 lln=1 lmax=1e-005 lmin=1.2e-006 lnoff=5.4545454e-007 lpclm=8.1927273e-008 lpdiblc2=4.4675455e-010 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lu0=1.3568182e-009 lua1=1.0963636e-016 lua=2.5898182e-016 luc1=6.8727273e-018 luc=5.9935909e-017 lvoffcv=-2.1818182e-007 lvth0=-4.0909091e-009 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=1.9454546 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.34150727 pdiblc1=0.1484 pdiblc2=7.8434545e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.010844318 ua1=1.4086364e-009 ua=6.2990182e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.4527273e-011 uc=-1.6606591e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0.021818182 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_14' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.model pmos_3p3.15 pmos a0=1.1534 a1=0 a2=0.99 acde=1 acnqsmod=0 agidl=1.5908e-011 ags=0.17736 alpha0=0.0018936 alpha1=0 at=12000 b0=0 b1=0 beta0=43.599 bgidl=1.3902e+009 binunit=2 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cf=0 cgbo=1e-013 cgdl=4e-011 cgdo=1.24e-010 cgidl=7.5 cgsl=4e-011 cgso=1.24e-010 cit=0 cjs=0.00094344 cjswgs=4.794e-010 cjsws=1.5078e-010 ckappad=0.6 ckappas=0.6 clc=1e-007 cle=0.6 delta=0.01 diomod=1 dlc=-8e-009 dlcig=1.5e-007 dmcg=1.5e-007 drout=0.56 dsub=0.3659 dvt0=2.8985 dvt0w=0 dvt1=0.23999 dvt1w=5300000 dvt2=-0.016 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1.12 egidl=0.1009 em=4.1e+007 epsrox=3.9 eta0=0.2541 etab=-0.15284 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=1.653e-007 jswgs=0 jsws=2.1207e-013 jtss=1e-011 jtsswgs=1e-011 jtssws=1e-011 k1=1.0069 k2=-0.035251 k3=0 k3b=0 keta=-0.0091505 kt1=-0.29993 kt1l=0 kt2=-0.013066 ku0=0 kvsat=0 kvth0=0 level=54 lint=0 ll=0 lln=1 lmax=5.0001e-005 lmin=1e-005 lpe0=3.2493e-008 lpeb=0 ltvoff=0 lw=0 lwl=0 lwn=1 minv=-0.1 mjs=0.32084 mjswgs=0.21964 mjsws=0.05 mobmod=0 moin=15 ndep=5.6e+017 nfactor=0.8 ngate=6e+019 njs=1 njts=20 njtssw=20 njtsswg=20 noff=2 noia='pmos_3p3_noia' noib='pmos_3p3_noib' noic='pmos_3p3_noic' nsd=1e+020 ntnoi=1 paramchk=1 pbs=0.69939 pbswgs=0.65 pbsws=0.8022 pclm=0.3497 pdiblc1=0.1484 pdiblc2=0.00012311 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0 prt=0 prwb=0 prwg=0 pscbe1=6.7448e+008 pscbe2=1e-005 ptvoff=0 pvag=0 rbodymod=0 rdsmod=0 rdsw='pmos_3p3_rdsw' rdswmin=20 rgatemod=0 rsh=7 saref=4.4e-007 sbref=4.4e-007 tcj=0.00099187 tcjsw=0.00063483 tcjswg=0.000932 tnoimod=0 tnom=25 toxe='pmos_3p3_tox' toxm=7.9e-009 toxp='pmos_3p3_tox' toxref=7.9e-009 tpb=0.0016906 tpbsw=0.0052 tpbswg=0.000744 trnqsmod=0 tvoff=0.0032 u0=0.01098 ua1=1.4196e-009 ua=6.558e-010 ub1=-2.6523e-018 ub=9.7125e-019 uc1=-6.384e-011 uc=-1.0613e-011 ute=-1 vbm=-3 version=4.5 vfb=0 vfbcv=-1 voff=-0.097861 voffcv=0 voffl=0 vsat=94000 vth0='pmos_3p3_vth0_15' vtss=10 vtsswgs=10 vtssws=10 w0=2.5e-006 wint=-1e-008 wl=0 wln=1 wmax=0.000100001 wmin=1e-005 wtvoff=0 ww=0 wwl=0 wwn=1 xj='pmos_3p3_xj' xl='pmos_3p3_xl' xpart=0 xtis=3 xw='pmos_3p3_xw'
.subckt pplus_u_m1 1 2 3 r_length='lr' r_width='wr' dtemp=0 par=1 r_rsh0='rsh_pplus_u_m' r_dw=2.75e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.375e-3 r_tc2=1e-6 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model pn_junction d cj=0.00094344 level=2
d1 1 3 pn_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends pplus_u_m1
.endl pmos_3p3_stat

.lib nmos_6p0_nat_stat
.subckt nmos_6p0_nat d g s b w=1e-5 l=1.8e-6 as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 par=1 dtemp=0 sa=0 sb=0 nf=1 sd=0 m=1
m0 d g s b nmos_6p0_nat m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' sa='sa' sb='sb' nf='nf' sd='sd'
.ends nmos_6p0_nat
.model nmos_6p0_nat.0 nmos a0=0.88 a1=0 a2=0.47 acde=0.3 acnqsmod=0 agidl=2e-010 ags=0.72 aigbacc=0.43 aigbinv=0.35 aigc=0.43 aigsd=0.43 alpha0=1.36e-008 alpha1=1e-005 at=80000 b0=3.5e-007 b1=0 beta0=15 bgidl=2.3e+009 bigbacc=0.054 bigbinv=0.03 bigc=0.054 bigsd=0.054 binunit=1 bvs=11 capmod=2 cdsc=0.00024 cdscb=0 cdscd=0 cgbo=1e-013 cgdl=1.5e-010 cgdo=1e-010 cgidl=0.5 cgsl=1.5e-010 cgso=1e-010 cigbacc=0.075 cigbinv=0.006 cigc=0.075 cigsd=0.075 cit=0 cjs=0.00095 cjswgs=3.573e-010 cjsws=1.33e-010 ckappad=0.6 ckappas=0.6 clc=1e-010 cle=0.6 delta=0.005 diomod=1 dlc=0 dlcig=0 dmcg=0 dmcgt=0 dmdg=0 drout=0.16 dsub=0.4 dvt0=2.2 dvt0w=0 dvt1=0.53 dvt1w=5300000 dvt2=-0.032 dvt2w=-0.032 dvtp0=1e-008 dvtp1=0 dwb=0 dwc=0 dwg=0 ef=1 egidl=0.8 eigbinv=1.1 em=4.1e+007 epsrox=3.9 eta0=0.06 etab=-0.43 eu=1.67 fnoimod=1 fprout=65 gbmin=1e-012 geomod=0 igbmod=0 igcmod=0 ijthsfwd=0.1 ijthsrev=0.1 jss=6.88e-007 jswgs=0 jsws=4.88e-013 jtsd=0 jtss=0 jtsswd=0 jtsswgd=0 jtsswgs=0 jtssws=0 k1=0.165 k2=-0.001 k2we=0 k3=-0.6 k3b=-0.6 keta=-0.04 kt1=-0.412 kt1l=3.5e-008 kt2=-0.05 ku0=0 ku0we=0 kvsat=0 kvth0=0 kvth0we=0 lambda=0 lat=-30000 level=54 lint=1e-007 lintnoi=0 lku0=0 lkvth0=0 ll=0 llc=0 lln=1 llodku0=0 llodvth=0 lmax=50.01e-6 lmin=1.8e-6 lnfactor=0.45 lodeta0=1 lodk2=1 lp=1e-008 lpe0=1e-007 lpeb=0 lu0=0.042 lub=3.65e-018 lute=-0.26 lvth0=-0.088 lw=0 lwc=0 lwl=0 lwlc=0 lwn=1 minv=-0.5 mjs=0.296 mjswgs=0.40313 mjsws=0.01 mobmod=0 moin=15 ndep=1.7e+017 nfactor=0.40241 ngate=1e+020 ngcon=1 nigbacc=1 nigbinv=3 nigc=1 njs=1.0541 njts=20 njtssw=20 njtsswg=20 noff=1.5 noia='nmos_6p0_nat_noia' noib='nmos_6p0_nat_noib' noic='nmos_6p0_nat_noic' nsd=1e+020 ntnoi=1 ntox=1 paramchk=1 pat=-10000 pbs=0.606 pbswgs=0.861 pbsws=0.48 pclm=3 pdiblc1=1.41 pdiblc2=1e-005 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 permod=1 phin=0.5 pigcd=1 pku0=0 pkvth0=0 poxedge=1 prt=0 prwb=0 prwg=1 pscbe1=5e+009 pscbe2=5e-006 pvag=1 pvsat=23500 rbdb=50 rbdbx0=100 rbdby0=100 rbodymod=0 rbpb=50 rbpbx0=100 rbpbxl=0 rbpbxnf=0 rbpbxw=0 rbpby0=100 rbpbyl=0 rbpbynf=0 rbpbyw=0 rbpd0=50 rbpd=50 rbpdl=0 rbpdnf=0 rbpdw=0 rbps0=50 rbps=50 rbpsl=0 rbpsnf=0 rbpsw=0 rbsb=50 rbsbx0=100 rbsby0=100 rbsdbxl=0 rbsdbxnf=0 rbsdbxw=0 rbsdbyl=0 rbsdbynf=0 rbsdbyw=0 rdsmod=0 rdsw='nmos_6p0_nat_rdsw' rdswmin=0 rdw=100 rdwmin=0 rgatemod=0 rsh=7 rshg=0.1 rsw=100 rswmin=0 saref=1e-006 sbref=1e-006 scref=1e-006 steta0=0 stk2=0 tcj=0.000825 tcjsw=0.0018 tcjswg=0.001595 tempmod=0 tku0=0 tnjts=0 tnjtssw=0 tnjtsswg=0 tnoimod=0 tnom=25 toxe='nmos_6p0_nat_tox' toxm=1.52e-008 toxp='8e-10+nmos_6p0_nat_tox' toxref=1.52e-008 tpb=0.00146 tpbsw=0.00313 tpbswg=0.0016588 trnqsmod=0 tvfbsdoff=0 tvoff=0 u0=0.070102 ua1=1e-009 ua=2.278e-009 ub1=-1e-018 ub=3.97e-019 uc1=-5.6e-011 uc=2.625e-012 ud1=0 up=0 ute=-1.5 vbm=-3 version=4.5 vfbcv=-1 vfbsdoff=0 voff=-0.06 voffcv=0 voffl=0 vsat=106700 vth0='nmos_6p0_nat_vth0' vtl=200000 vtsd=10 vtss=10 vtsswd=10 vtsswgd=10 vtsswgs=10 vtssws=10 w0=1e-010 web=0 wec=0 wint=1e-009 wku0=0 wkvth0=0 wl=0 wlc=0 wln=1 wlod=0 wlodku0=0 wlodvth=0 wmax=100.01e-6 wmin=0.8e-6 wpemod=0 wr=1 ww=0 wwc=0 wwl=0 wwlc=0 wwn=1 xgl=0 xgw=0 xj='nmos_6p0_nat_xj' xjbvd=1 xjbvs=1 xl='nmos_6p0_nat_xl' xn=3 xpart=0 xrcrg1=12 xrcrg2=1 xtis=3 xtsd=0.02 xtss=0.02 xtsswd=0.02 xtsswgd=0.02 xtsswgs=0.02 xtssws=0.02 xw='nmos_6p0_nat_xw'
.endl nmos_6p0_nat_stat

.lib pmos_6p0_stat
.subckt pmos_6p0_sab d g s b w=10u l=0.5u par=1 s_sab=0.28u d_sab=2.78u as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 dtemp=0 nf=1 sa=0 sb=0 sd=0 m=1
.param par_vth=0.01051
.param par_k=0.00517
.param par_l=3e-7
.param par_w=-4e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
xr1 d d1 b pplus_u_m2 wr='w' lr='(d_sab==0)?1e-15:d_sab' dtemp='dtemp'
xr2 s s1 b pplus_u_m2 wr='w' lr='(s_sab==0)?1e-15:s_sab' dtemp='dtemp'
m0 d1 g s1 b pmos_6p0 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' nf='nf' sa='0' sb='0' sd='0' delvto='mis_vth*sw_stat_mismatch'
.ends
.model pmos_6p0.0 pmos a0=0.84 a1=0 a2=1 acde=0.7 acnqsmod=0 ags=0.059 alpha0=9.6e-7 alpha1=51.5 at=-2.18e4 b0=2.625e-8 b1=0 beta0=50.8 binunit=1 bvd=10.5 bvs=10.5 capmod=2 cdsc=2.4e-4 cdscb=0 cdscd=0 cgbo=1e-13 cgdl=5.25e-11 cgdo=7.71e-11 cgsl=5.25e-11 cgso=7.71e-11 cit=0 cjd=0.000912 cjs=0.000912 cjswd=1.4649e-010 cjswgd=3.3229e-010 cjswgs=3.3229e-010 cjsws=1.4649e-010 ckappad=0.6 ckappas=0.6 delta=0.01 diomod=1 dlc=7.4e-9 drout=0.56 dsub=0.4824 dvt0=1 dvt0w=0 dvt1=1 dvt1w=5.3e6 dvt2=0 dvt2w=-0.032 dvtp0=0 dvtp1=0.3 dwb=-3e-9 dwg=-6.6e-9 ef=1.1 epsrox=3.9 eta0=0.08 etab=-0.09408 fnoimod=1 fprout=0 geomod=1 igbmod=0 igcmod=0 ijthdfwd=0.1 ijthdrev=0.1 ijthsfwd=0.1 ijthsrev=0.1 jsd=2.0867e-007 jss=2.0867e-007 jswd=1.6088e-013 jswgd=0 jswgs=0 jsws=1.6088e-013 k1=0.9588 k2=8.936e-3 k3=-0.75 k3b=1.2104 keta=-8.6016e-5 kt1=-0.3828 kt1l=-3.158e-8 kt2=-0.09064 lambda=0 lc=0 level=54 lint=6.7e-8 ll=-5.4e-15 lln=1 lmax=50.01e-6 lmin=0.5e-6 lpe0=-4.4e-8 lpeb=-5.96e-8 lphin=0.1408 lua1=-6.554813e-10 lub1=1.939773e-19 luc1=-1.067674e-10 luc=8.691408e-11 lute=-0.152467 lw=0 lwl=-4.76e-21 lwn=1 minv=0 mjd=0.32713 mjs=0.32713 mjswd=0.056777 mjswgd=0.50996 mjswgs=0.50996 mjsws=0.056777 mobmod=0 moin=15 ndep=1.7e17 nfactor=1 ngate=3.6e19 njd=1 njs=1 noff=1 noia='pmos_6p0_noia' noib='pmos_6p0_noib' noic='pmos_6p0_noic' nsd=6e16 paramchk=1 pat=-6.1e3 pbd=0.76836 pbeta0=0.14 pbs=0.76836 pbswd=0.5 pbswgd=1.2295 pbswgs=1.2295 pbsws=0.5 pclm=0.42 pdiblc1=0.14 pdiblc2=1e-5 pdiblcb=0 pdits=0.01 pditsd=0 pditsl=0 permod=1 petab=-0.012128 phin=0 pkt1=2.2e-3 ppclm=0.071 pprwb=-0.052 prdsw=-120 prt=454 prwb=0.569552 prwg=0.0432 pscbe1=5.088e8 pscbe2=1e-8 pua1=-3.823641e-10 pub1=7.291324e-19 puc1=1.8536e-11 puc=-1.501336e-11 pvag=1.5 pvth0=7.6e-3 rbodymod=0 rdsmod=0 rdsw='pmos_6p0_rdsw' rdswmin=100 rsh=7 rshg=0.1 tcj=0.001 tcjsw=0.00071888 tcjswg=0.0009411 tempmod=0 tnoimod=0 tnom=25 toxe='pmos_6p0_tox' tpb=0.0019314 tpbsw=0.0017642 tpbswg=0.0016588 trnqsmod=0 u0=0.0151 ua1=1.41e-9 ua=1.78e-9 ub1=-4.31e-18 ub=4.88e-19 uc1=1.147552e-10 uc=-2.7435e-11 ute=-1.2 version=4.5 vfb=-1 voff=-0.1284 voffcv=0 voffl=2.19e-8 vsat=8.55e4 vth0='pmos_6p0_vth0' vtl=2e5 w0=3.1e-7 wbeta0=0.22 wint=4.9e-8 wketa=2.772e-3 wl=0 wln=1 wmax=100.01e-6 wmin=0.3e-6 wr=1 wrdsw=213.9 wua1=-1.2e-10 wute=-0.07 ww=-1.37e-14 wwl=3.04e-22 wwn=1 xj='pmos_6p0_xj' xjbvd=1 xjbvs=1 xl='pmos_6p0_xl' xn=3 xpart=1 xtid=3 xtis=3 xw='pmos_6p0_xw'
.subckt pplus_u_m2 1 2 3 r_length='lr' r_width='wr' dtemp=0 par=1 r_rsh0='rsh_pplus_u_m' r_dw=2.75e-8 r_dl=0 r_vc1=0 r_vc2=0 r_tc1=1.375e-3 r_tc2=1e-6 r_tnom=25 r_l='r_length-2*r_dl' r_w='r_width-2*r_dw' r_n='r_l/r_w' r_temp='1+r_tc1*(temp+dtemp-r_tnom)+r_tc2*(temp+dtemp-r_tnom)*(temp+dtemp-r_tnom)'
.model pn_junction d cj=0.00094344 level=2
d1 1 3 pn_junction area='r_w*r_l'
rb 1 2 r='r_temp*r_n*(r_rsh0+r_vc1*abs(v(1,2))/r_n+r_vc2*abs(v(1,2))*abs(v(1,2))/r_n/r_n)'
.ends pplus_u_m2
.endl pmos_6p0_stat

.lib efuse
.subckt efuse in out pblow=0
rfuse in out r='200*(1-pblow)+900*pblow'
.ends efuse
.endl efuse

.lib fets_mm
.subckt nmos_3p3 d g s b w=1e-5 l=2.8e-7 as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 par=1 dtemp=0 sa=0 sb=0 nf=1 sd=0 m=1
.param par_vth=0.007148
.param par_k=0.007008
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
m0 d g s b nmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' delvto='mis_vth*sw_stat_mismatch' sa='sa' sb='sb' nf='nf' sd='sd'
.ends nmos_3p3
.subckt pmos_3p3 d g s b w=1e-5 l=2.8e-7 as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 par=1 dtemp=0 sa=0 sb=0 nf=1 sd=0 m=1
.param par_vth=0.00666
.param par_k=0.002833
.param par_l=1.5e-7
.param par_w=-1e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
m0 d g s b pmos_3p3 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' delvto='mis_vth*sw_stat_mismatch' sa='sa' sb='sb' nf='nf' sd='sd'
.ends pmos_3p3
.subckt nmos_6p0 d g s b w=1e-5 l=7e-7 as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 par=1 dtemp=0 sa=0 sb=0 nf=1 sd=0 m=1
.param par_vth=0.01155
.param par_k=0.0000
.param par_l=4e-7
.param par_w=-5e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
m0 d g s b nmos_6p0 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' delvto='mis_vth*sw_stat_mismatch' sa='sa' sb='sb' nf='nf' sd='sd'
.ends nmos_6p0
.subckt pmos_6p0 d g s b w=1e-5 l=5e-7 as=0 ad=0 ps=0 pd=0 nrd=0 nrs=0 par=1 dtemp=0 sa=0 sb=0 nf=1 sd=0 m=1
.param par_vth=0.01051
.param par_k=0.00517
.param par_l=3e-7
.param par_w=-4e-7
.param par_leff='l-par_l'
.param par_weff='par*(w-par_w)'
.param p_sqrtarea='sqrt((par_leff)*(par_weff))'
.param var_k='0.7071*par_k*1e-06/p_sqrtarea'
.param mis_k='agauss(0,var_k,1)'
.param var_vth='0.7071*par_vth*1e-06/p_sqrtarea'
.param mis_vth='agauss(0,var_vth,1)'
m0 d g s b pmos_6p0 m='m' w='w' l='l' as='as' ad='ad' ps='ps' pd='pd' nrd='nrd' nrs='nrs' delvto='mis_vth*sw_stat_mismatch' sa='sa' sb='sb' nf='nf' sd='sd'
.ends pmos_6p0
.endl fets_mm

.lib res_statistical_par
.param mc_rsh_nplus_u=0
.param mc_rsh_pplus_u=0
.param mc_rsh_nplus_s=0
.param mc_rsh_pplus_s=0
.param mc_rsh_npolyf_u=0
.param mc_rsh_ppolyf_u=0
.param mc_rsh_npolyf_s=0
.param mc_rsh_ppolyf_s=0
.param mc_rsh_ppolyf_u_1k=0
.param mc_rsh_ppolyf_u_2k=0
.param mc_rsh_ppolyf_u_1k_6p0=0
.param mc_rsh_ppolyf_u_2k_6p0=0
.param mc_rsh_ppolyf_u_3k=0
.param mc_dw_nplus_u=0
.param mc_dw_pplus_u=0
.param mc_dw_nplus_s=0
.param mc_dw_pplus_s=0
.param mc_dw_npolyf_u=0
.param mc_dw_ppolyf_u=0
.param mc_dw_npolyf_s=0
.param mc_dw_ppolyf_s=0
.param mc_dw_ppolyf_u_1k=0
.param mc_dw_ppolyf_u_2k=0
.param mc_dw_ppolyf_u_1k_6p0=0
.param mc_dw_ppolyf_u_2k_6p0=0
.param mc_dw_ppolyf_u_3k=0
.param mc_rt_nplus_u=0
.param mc_rt_pplus_u=0
.param mc_rt_npolyf_u=0
.param mc_rt_ppolyf_u=0
.param mc_rt_ppolyf_u_1k=0
.param mc_rt_ppolyf_u_2k=0
.param mc_rt_ppolyf_u_1k_6p0=0
.param mc_rt_ppolyf_u_2k_6p0=0
.param mc_rt_ppolyf_u_3k=0
.endl res_statistical_par

.lib res_statistical
.param rsh_nplus_u=60
.param rsh_pplus_u=185
.param rsh_nplus_s=6.3
.param rsh_pplus_s=7
.param rsh_nwell=1000
.param rsh_npolyf_u=310
.param rsh_ppolyf_u=350
.param rsh_npolyf_s=6.8
.param rsh_ppolyf_s=7.3
.param rsh_ppolyf_u_1k=1000
.param rsh_ppolyf_u_2k=2000
.param rsh_ppolyf_u_1k_6p0=1000
.param rsh_ppolyf_u_2k_6p0=2000
.param rsh_ppolyf_u_3k=3000
.param rsh_rm1=0.09
.param rsh_rm2=0.09
.param rsh_rm3=0.09
.param rsh_tm6k=60e-3
.param rsh_tm9k=40e-3
.param rsh_tm11k=40e-3
.param rsh_tm30k=9.5e-3
.param mc_rsh_nplus_u_temp='agauss(0,3.8,3)'
.param mc_rsh_pplus_u_temp='agauss(0,10.055,3)'
.param mc_rsh_nplus_s_temp='agauss(0,1.33,3)'
.param mc_rsh_pplus_s_temp='agauss(0,1.4917,3)'
.param mc_rsh_npolyf_u_temp='agauss(0,15.135,3)'
.param mc_rsh_ppolyf_u_temp='agauss(0,18.116,3)'
.param mc_rsh_npolyf_s_temp='agauss(0,1.392,3)'
.param mc_rsh_ppolyf_s_temp='agauss(0,1.5852,3)'
.param mc_rsh_ppolyf_u_1k_temp='agauss(0,49.754,3)'
.param mc_rsh_ppolyf_u_2k_temp='agauss(0,101.518,3)'
.param mc_rsh_ppolyf_u_1k_6p0_temp='agauss(0,51.894,3)'
.param mc_rsh_ppolyf_u_2k_6p0_temp='agauss(0,99.242,3)'
.param mc_rsh_ppolyf_u_3k_temp='agauss(0,184.603,3)'
.param mc_dw_nplus_u_temp='agauss(0,0.0144,3)'
.param mc_dw_pplus_u_temp='agauss(0,0.0144,3)'
.param mc_dw_nplus_s_temp='agauss(0,0.012,3)'
.param mc_dw_pplus_s_temp='agauss(0,0.018,3)'
.param mc_dw_npolyf_u_temp='agauss(0,0.0167,3)'
.param mc_dw_ppolyf_u_temp='agauss(0,0.0167,3)'
.param mc_dw_npolyf_s_temp='agauss(0,0.006,3)'
.param mc_dw_ppolyf_s_temp='agauss(0,0.003,3)'
.param mc_dw_ppolyf_u_1k_temp='agauss(0,0.0167,3)'
.param mc_dw_ppolyf_u_2k_temp='agauss(0,0.0167,3)'
.param mc_dw_ppolyf_u_1k_6p0_temp='agauss(0,0.0167,3)'
.param mc_dw_ppolyf_u_2k_6p0_temp='agauss(0,0.0167,3)'
.param mc_dw_ppolyf_u_3k_temp='agauss(0,0.0167,3)'
.param mc_rt_nplus_u_temp='agauss(0,0.64,3)'
.param mc_rt_pplus_u_temp='agauss(0,7.2,3)'
.param mc_rt_npolyf_u_temp='agauss(0,4.8,3)'
.param mc_rt_ppolyf_u_temp='agauss(0,4.7,3)'
.param mc_rt_ppolyf_u_1k_temp='agauss(0,6.838,3)'
.param mc_rt_ppolyf_u_2k_temp='agauss(0,6.838,3)'
.param mc_rt_ppolyf_u_1k_6p0_temp='agauss(0,6.838,3)'
.param mc_rt_ppolyf_u_2k_6p0_temp='agauss(0,6.838,3)'
.param mc_rt_ppolyf_u_3k_temp='agauss(0,6.93,3)'
.param mc_rsh_nplus_u='mc_rsh_nplus_u_temp'
.param mc_rsh_pplus_u='mc_rsh_pplus_u_temp'
.param mc_rsh_nplus_s='mc_rsh_nplus_s_temp'
.param mc_rsh_pplus_s='mc_rsh_pplus_s_temp'
.param mc_rsh_npolyf_u='mc_rsh_npolyf_u_temp'
.param mc_rsh_ppolyf_u='mc_rsh_ppolyf_u_temp'
.param mc_rsh_npolyf_s='mc_rsh_npolyf_s_temp'
.param mc_rsh_ppolyf_s='mc_rsh_ppolyf_s_temp'
.param mc_rsh_ppolyf_u_1k='mc_rsh_ppolyf_u_1k_temp'
.param mc_rsh_ppolyf_u_2k='mc_rsh_ppolyf_u_2k_temp'
.param mc_rsh_ppolyf_u_1k_6p0='mc_rsh_ppolyf_u_1k_6p0_temp'
.param mc_rsh_ppolyf_u_2k_6p0='mc_rsh_ppolyf_u_2k_6p0_temp'
.param mc_rsh_ppolyf_u_3k='mc_rsh_ppolyf_u_3k_temp'
.param mc_dw_nplus_u='mc_dw_nplus_u_temp'
.param mc_dw_pplus_u='mc_dw_pplus_u_temp'
.param mc_dw_nplus_s='mc_dw_nplus_s_temp'
.param mc_dw_pplus_s='mc_dw_pplus_s_temp'
.param mc_dw_npolyf_u='mc_dw_npolyf_u_temp'
.param mc_dw_ppolyf_u='mc_dw_ppolyf_u_temp'
.param mc_dw_npolyf_s='mc_dw_npolyf_s_temp'
.param mc_dw_ppolyf_s='mc_dw_ppolyf_s_temp'
.param mc_dw_ppolyf_u_1k='mc_dw_ppolyf_u_1k_temp'
.param mc_dw_ppolyf_u_2k='mc_dw_ppolyf_u_2k_temp'
.param mc_dw_ppolyf_u_1k_6p0='mc_dw_ppolyf_u_1k_6p0_temp'
.param mc_dw_ppolyf_u_2k_6p0='mc_dw_ppolyf_u_2k_6p0_temp'
.param mc_dw_ppolyf_u_3k='mc_dw_ppolyf_u_3k_temp'
.param mc_rt_nplus_u='mc_rt_nplus_u_temp'
.param mc_rt_pplus_u='mc_rt_pplus_u_temp'
.param mc_rt_npolyf_u='mc_rt_npolyf_u_temp'
.param mc_rt_ppolyf_u='mc_rt_ppolyf_u_temp'
.param mc_rt_ppolyf_u_1k='mc_rt_ppolyf_u_1k_temp'
.param mc_rt_ppolyf_u_2k='mc_rt_ppolyf_u_2k_temp'
.param mc_rt_ppolyf_u_1k_6p0='mc_rt_ppolyf_u_1k_6p0_temp'
.param mc_rt_ppolyf_u_2k_6p0='mc_rt_ppolyf_u_2k_6p0_temp'
.param mc_rt_ppolyf_u_3k='mc_rt_ppolyf_u_3k_temp'
.lib 'sm141064.spice' res
.lib 'sm141064.spice' efuse
.endl res_statistical

.lib bjt_statistical
.param isa=1
.param bfa=1
.param rba=1
.param rea=1
.param rca=1
.param rbma=1
.param cjea=1
.param cjca=1
.param is_cor_npn=1
.param bf_cor_npn=1
.param rb_cor_npn=1
.param re_cor_npn=1
.param rc_cor_npn=1
.param rbm_cor_npn=1
.param cjc_cor_npn=1
.param cje_cor_npn=1
.param mc_xis_vnpn_temp='agauss(0,0.7,3)'
.param mc_xbf_vnpn_temp='agauss(0,0.48,3)'
.param mc_xrb_vnpn_temp='agauss(0,0.2,3)'
.param mc_xre_vnpn_temp='agauss(0,0.2,3)'
.param mc_xrc_vnpn_temp='agauss(0,0.2,3)'
.param mc_xcje_vnpn_temp='agauss(0,0.15,3)'
.param mc_xcjc_vnpn_temp='agauss(0,0.15,3)'
.param mc_xis_vpnp_temp='agauss(0,0.3,3)'
.param mc_xbf_vpnp_temp='agauss(0,0.2,3)'
.param mc_xrb_vpnp_temp='agauss(0,0.2,3)'
.param mc_xre_vpnp_temp='agauss(0,0.2,3)'
.param mc_xrc_vpnp_temp='agauss(0,0.2,3)'
.param mc_xcje_vpnp_temp='agauss(0,0.15,3)'
.param mc_xcjc_vpnp_temp='agauss(0,0.15,3)'
.param mc_xis_vnpn='mc_xis_vnpn_temp'
.param mc_xbf_vnpn='mc_xbf_vnpn_temp'
.param mc_xrb_vnpn='mc_xrb_vnpn_temp'
.param mc_xre_vnpn='mc_xre_vnpn_temp'
.param mc_xrc_vnpn='mc_xrc_vnpn_temp'
.param mc_xcje_vnpn='mc_xcje_vnpn_temp'
.param mc_xcjc_vnpn='mc_xcjc_vnpn_temp'
.param mc_xis_vpnp='mc_xis_vpnp_temp'
.param mc_xbf_vpnp='mc_xbf_vpnp_temp'
.param mc_xrb_vpnp='mc_xrb_vpnp_temp'
.param mc_xre_vpnp='mc_xre_vpnp_temp'
.param mc_xrc_vpnp='mc_xrc_vpnp_temp'
.param mc_xcje_vpnp='mc_xcje_vpnp_temp'
.param mc_xcjc_vpnp='mc_xcjc_vpnp_temp'
.lib 'sm141064.spice' bjt_mc
.endl bjt_statistical

.lib bjt_mc
.subckt vpnp_0p42x10 c b e par=1 dtemp=0
.param mis_is_vpnp_0p42x10='agauss(0,0.0015,1)'
.param mis_bf_vpnp_0p42x10='agauss(0,0.01088,1)'
.param isa_mis_vpnp_0p42x10='mis_is_vpnp_0p42x10*sw_stat_mismatch/sqrt(par)'
.param bf_mis_vpnp_0p42x10='mis_bf_vpnp_0p42x10*sw_stat_mismatch/sqrt(par)'
q0 c b e vpnp_0p42x10
.model vpnp_0p42x10 pnp af=1 bf='1.69*bfa*(1+mc_xbf_vpnp*sw_stat_global)*(1+bf_mis_vpnp_0p42x10)' br=0.0036 cjc='2.04e-014*cjca*(1+mc_xcjc_vpnp*sw_stat_global)' cje='6.88e-015*cjea*(1+mc_xcje_vpnp*sw_stat_global)' cjs=0 eg=1.17 fc=0.5 ikf=0.00063375 ikr=0.1 irb=0.1 is='9e-019*isa*(1+mc_xis_vpnp*sw_stat_global)*(1+isa_mis_vpnp_0p42x10)' isc=1e-018 ise=2.7e-016 itf=0.1 kf=0 mjc=0.22711 mje=0.14469 mjs=0.5 nc=2 ne=1.64 nf=1 nkf=0.4 nr=1 ptf=0 rb='41*rba*(1+mc_xrb_vpnp*sw_stat_global)' rbm='10*rbma' rc='10*rca*(1+mc_xrc_vpnp*sw_stat_global)' re='1*rea*(1+mc_xre_vpnp*sw_stat_global)' tf=1e-010 tr=0 vaf=80 var=23 vjc=0.43905 vje=0.43905 vjs=0.75 vtf=10 xcjc=1 xtb=0.0001 xtf=1 xti=3 level=1
.ends vpnp_0p42x10
.subckt vpnp_0p42x5 c b e par=1 dtemp=0
.param mis_is_vpnp_0p42x5='agauss(0,0.0017,1)'
.param mis_bf_vpnp_0p42x5='agauss(0,0.0119,1)'
q0 c b e vpnp_0p42x5
.model vpnp_0p42x5 pnp af=1 bf='1.681*bfa*(1+mc_xbf_vpnp*sw_stat_global)*(1+mis_bf_vpnp_0p42x5*sw_stat_mismatch/sqrt(par))' br=1.9872e-3 cjc='1.17e-14*cjca*(1+mc_xcjc_vpnp*sw_stat_global)' cje='3.5e-15*cjea*(1+mc_xcje_vpnp*sw_stat_global)' cjs=0 eg=1.17 fc=0.5 ikf=2.4777e-4 ikr=0.1 irb=0.1 is='4.388e-19*isa*(1+mc_xis_vpnp*sw_stat_global)*(1+mis_is_vpnp_0p42x5*sw_stat_mismatch/sqrt(par))' isc=1e-16 ise=1.2124e-16 itf=0.1 kf=0 mjc=0.22711 mje=0.15395 mjs=0.5 nc=2 ne=1.64 nf=1 nkf=0.4 nr=1 ptf=0 rb='41*rba*(1+mc_xrb_vpnp*sw_stat_global)' rbm='10*rbma' rc='10*rca*(1+mc_xrc_vpnp*sw_stat_global)' re='1*rea*(1+mc_xre_vpnp*sw_stat_global)' tf=1e-10 tr=0 vaf=180 var=23 vjc=0.43905 vje=0.43905 vjs=0.75 vtf=10 xcjc=1 xtb=1e-4 xtf=1 xti=3 level=1
.ends vpnp_0p42x5
.subckt vpnp_10x10 c b e par=1 dtemp=0
.param mis_is_vpnp_10x10='agauss(0,0.00077,1)'
.param mis_bf_vpnp_10x10='agauss(0,0.0013,1)'
q0 c b e vpnp_10x10
.model vpnp_10x10 pnp af=1 bf='1.7*bfa*(1+mc_xbf_vpnp*sw_stat_global)*(1+mis_bf_vpnp_10x10*sw_stat_mismatch/sqrt(par))' br=0.017038 cjc='4.69e-14*cjca*(1+mc_xcjc_vpnp*sw_stat_global)' cje='9.71e-14*cjea*(1+mc_xcje_vpnp*sw_stat_global)' cjs=0 eg=1.17 fc=0.5 ikf=2.610625e-3 ikr=0.1 irb=0.1 is='1.249175e-17*isa*(1+mc_xis_vpnp*sw_stat_global)*(1+mis_is_vpnp_10x10*sw_stat_mismatch/sqrt(par))' isc=1e-18 ise=2.7e-16 itf=0.1 kf=0 mjc=0.24528 mje=0.24192 mjs=0.5 nc=2 ne=1.64 nf=1 nkf=0.4 nr=1 ptf=0 rb='27.88*rba*(1+mc_xrb_vpnp*sw_stat_global)' rbm='10*rbma' rc='10*rca*(1+mc_xrc_vpnp*sw_stat_global)' re='1*rea*(1+mc_xre_vpnp*sw_stat_global)' tf=1e-10 tr=0 vaf=206.4 var=23 vjc=0.43905 vje=0.43905 vjs=0.75 vtf=10 xcjc=1 xtb=1e-4 xtf=1 xti=3 level=1
.ends vpnp_10x10
.subckt vpnp_5x5 c b e par=1 dtemp=0
.param mis_is_vpnp_5x5='agauss(0,0.00052,1)'
.param mis_bf_vpnp_5x5='agauss(0,0.0031,1)'
q0 c b e vpnp_5x5
.model vpnp_5x5 pnp af=1 bf='1.65*bfa*(1+mc_xbf_vpnp*sw_stat_global)*(1+mis_bf_vpnp_5x5*sw_stat_mismatch/sqrt(par))' br=8.372e-3 cjc='2.15e-14*cjca*(1+mc_xcjc_vpnp*sw_stat_global)' cje='2.57e-14*cjea*(1+mc_xcje_vpnp*sw_stat_global)' cjs=0 eg=1.17 fc=0.5 ikf=1.025275e-3 ikr=0.1 irb=0.1 is='3.403e-18*isa*(1+mc_xis_vpnp*sw_stat_global)*(1+mis_is_vpnp_5x5*sw_stat_mismatch/sqrt(par))' isc=1e-18 ise=2.7e-16 itf=0.1 kf=0 mjc=0.22711 mje=0.23266 mjs=0.5 nc=2 ne=1.64 nf=1 nkf=0.4 nr=1 ptf=0 rb='41*rba*(1+mc_xrb_vpnp*sw_stat_global)' rbm='10*rbma' rc='10*rca*(1+mc_xrc_vpnp*sw_stat_global)' re='1*rea*(1+mc_xre_vpnp*sw_stat_global)' tf=1e-10 tr=0 vaf=208.8 var=27.37 vjc=0.43905 vje=0.43905 vjs=0.75 vtf=10 xcjc=1 xtb=1e-4 xtf=1 xti=3 level=1
.ends vpnp_5x5
.subckt vnpn_10x10 c b e s par=1 dtemp=0
q0 c b e s vnpn_10x10
.model vnpn_10x10 npn af=1 bf='10.83*bf_cor_npn*(1+mc_xbf_vnpn*sw_stat_global)' br=0.258 cjc='7.053e-14*cjc_cor_npn*(1+mc_xcjc_vnpn*sw_stat_global)' cje='1.031e-13*cje_cor_npn*(1+mc_xcje_vnpn*sw_stat_global)' cjs=1.135e-13 eg=1.17 ikf=0.021028 ikr=0.0038951 irb=0.00045303 is='1.8108e-017*is_cor_npn*(1+mc_xis_vnpn*sw_stat_global)' isc=1.5816e-016 ise=2.9626e-016 kf=0 mjc=0.31113 mje=0.32071 mjs=0.14716 nc=1.284 ne=1.345 nf=1.002 nkf=0.584 nr=1.002 rb='65.442*rb_cor_npn*(1+mc_xrb_vnpn*sw_stat_global)' rbm='1*rbm_cor_npn' rc='10.146*rc_cor_npn*(1+mc_xrc_vnpn*sw_stat_global)' re='6.9007*re_cor_npn*(1+mc_xre_vnpn*sw_stat_global)' vaf=95.696 var=29.681 vjc=0.63391 vje=0.70172 vjs=0.35175 xcjc=1 xtb=0 xti=3 level=1
.ends vnpn_10x10
.subckt vnpn_5x5 c b e s par=1 dtemp=0
q0 c b e s vnpn_5x5
.model vnpn_5x5 npn af=1 bf='10.05*bf_cor_npn*(1+mc_xbf_vnpn*sw_stat_global)' br=0.16573 cjc='2.972e-14*cjc_cor_npn*(1+mc_xcjc_vnpn*sw_stat_global)' cje='2.733e-14*cje_cor_npn*(1+mc_xcje_vnpn*sw_stat_global)' cjs=6.618e-14 eg=1.17 ikf=0.01158 ikr=0.0038951 irb=0.00045303 is='5.1456e-018*is_cor_npn*(1+mc_xis_vnpn*sw_stat_global)' isc=1.2536e-016 ise=2.5923e-016 kf=0 mjc=0.31113 mje=0.32071 mjs=0.14716 nc=1.284 ne=1.4224 nf=1.002 nkf=0.584 nr=1 rb='71.419*rb_cor_npn*(1+mc_xrb_vnpn*sw_stat_global)' rbm='1*rbm_cor_npn' rc='12.655*rc_cor_npn*(1+mc_xrc_vnpn*sw_stat_global)' re='12.809*re_cor_npn*(1+mc_xre_vnpn*sw_stat_global)' vaf=77.796 var=28.001 vjc=0.63391 vje=0.70172 vjs=0.35175 xcjc=1 xtb=0 xti=3 level=1
.ends vnpn_5x5
.subckt vnpn_0p54x16 c b e s par=1 dtemp=0
q0 c b e s vnpn_0p54x16
.model vnpn_0p54x16 npn af=1 bf='8.4987*bf_cor_npn*(1+mc_xbf_vnpn*sw_stat_global)' br=0.079582 cjc='3.540e-14*cjc_cor_npn*(1+mc_xcjc_vnpn*sw_stat_global)' cje='1.354e-14*cje_cor_npn*(1+mc_xcje_vnpn*sw_stat_global)' cjs=8.211e-14 eg=1.17 ikf=0.013121 ikr=0.0038951 irb=0.00045303 is='2.8872e-018*is_cor_npn*(1+mc_xis_vnpn*sw_stat_global)' isc=1.0425e-016 ise=5.2003e-016 kf=0 mjc=0.31113 mje=0.32071 mjs=0.14716 nc=1.284 ne=1.4678 nf=1.002 nkf=0.584 nr=1 rb='137.43*rb_cor_npn*(1+mc_xrb_vnpn*sw_stat_global)' rbm='1*rbm_cor_npn' rc='12.9*rc_cor_npn*(1+mc_xrc_vnpn*sw_stat_global)' re='14.121*re_cor_npn*(1+mc_xre_vnpn*sw_stat_global)' vaf=37.389 var=23.969 vjc=0.63391 vje=0.70172 vjs=0.35175 xcjc=1 xtb=0 xti=3 level=1
.ends vnpn_0p54x16
.subckt vnpn_0p54x8 c b e s par=1 dtemp=0
q0 c b e s vnpn_0p54x8
.model vnpn_0p54x8 npn af=1 bf='8.4*bf_cor_npn*(1+mc_xbf_vnpn*sw_stat_global)' br=0.069974 cjc='2.064e-14*cjc_cor_npn*(1+mc_xcjc_vnpn*sw_stat_global)' cje='6.857e-15*cje_cor_npn*(1+mc_xcje_vnpn*sw_stat_global)' cjs=5.703e-14 eg=1.17 ikf=0.0077487 ikr=0.0038951 irb=0.00045303 is='1.4309e-018*is_cor_npn*(1+mc_xis_vnpn*sw_stat_global)' isc=7.3712e-017 ise=2.6232e-016 kf=0 mjc=0.31113 mje=0.32071 mjs=0.14716 nc=1.284 ne=1.4685 nf=1.001 nkf=0.584 nr=0.996 rb='141.94*rb_cor_npn*(1+mc_xrb_vnpn*sw_stat_global)' rbm='1*rbm_cor_npn' rc='13.434*rc_cor_npn*(1+mc_xrc_vnpn*sw_stat_global)' re='14.573*re_cor_npn*(1+mc_xre_vnpn*sw_stat_global)' vaf=37.389 var=25.201 vjc=0.63391 vje=0.70172 vjs=0.35175 xcjc=1 xtb=0 xti=3 level=1
.ends vnpn_0p54x8
.subckt vnpn_0p54x4 c b e s par=1 dtemp=0
q0 c b e s vnpn_0p54x4
.model vnpn_0p54x4 npn af=1 bf='8.39*bf_cor_npn*(1+mc_xbf_vnpn*sw_stat_global)' br=0.057751 cjc='1.326e-14*cjc_cor_npn*(1+mc_xcjc_vnpn*sw_stat_global)' cje='3.513e-15*cje_cor_npn*(1+mc_xcje_vnpn*sw_stat_global)' cjs=4.449e-14 eg=1.17 ikf=0.0048817 ikr=0.0038951 irb=0.00045303 is='7.6696e-019*is_cor_npn*(1+mc_xis_vnpn*sw_stat_global)' isc=6.2655e-017 ise=1.3419e-016 kf=0 mjc=0.31113 mje=0.32071 mjs=0.14716 nc=1.284 ne=1.4801 nf=1.001 nkf=0.584 nr=0.998 rb='167*rb_cor_npn*(1+mc_xrb_vnpn*sw_stat_global)' rbm='1*rbm_cor_npn' rc='14.542*rc_cor_npn*(1+mc_xrc_vnpn*sw_stat_global)' re='17.058*re_cor_npn*(1+mc_xre_vnpn*sw_stat_global)' vaf=37.389 var=25.201 vjc=0.63391 vje=0.70172 vjs=0.35175 xcjc=1 xtb=0 xti=3 level=1
.ends vnpn_0p54x4
.subckt vnpn_0p54x2 c b e s par=1 dtemp=0
q0 c b e s vnpn_0p54x2
.model vnpn_0p54x2 npn af=1 bf='8.25*bf_cor_npn*(1+mc_xbf_vnpn*sw_stat_global)' br=0.043698 cjc='9.569e-15*cjc_cor_npn*(1+mc_xcjc_vnpn*sw_stat_global)' cje='1.841e-15*cje_cor_npn*(1+mc_xcje_vnpn*sw_stat_global)' cjs=3.822e-14 eg=1.17 ikf=0.0039054 ikr=0.0038951 irb=0.00045303 is='4.5765e-019*is_cor_npn*(1+mc_xis_vnpn*sw_stat_global)' isc=6.2655e-017 ise=8e-017 kf=0 mjc=0.31113 mje=0.32071 mjs=0.14716 nc=1.284 ne=1.49 nf=1.004 nkf=0.584 nr=1.0005 rb='231.74*rb_cor_npn*(1+mc_xrb_vnpn*sw_stat_global)' rbm='1*rbm_cor_npn' rc='17.312*rc_cor_npn*(1+mc_xrc_vnpn*sw_stat_global)' re='25.055*re_cor_npn*(1+mc_xre_vnpn*sw_stat_global)' vaf=37.389 var=25.201 vjc=0.63391 vje=0.70172 vjs=0.35175 xcjc=1 xtb=0 xti=3 level=1
.ends vnpn_0p54x2
.endl bjt_mc

.lib mimcap_statistical
.param mim_corner_1p5ff=1
.param mim_corner_1p0ff=1
.param mim_corner_2p0ff=1
.param mc_c_cox_1p0ff2='agauss(0,0.025,3)'
.param mc_c_cox_1p5ff2='agauss(0,0.03875,3)'
.param mc_c_cox_2p0ff2='agauss(0,0.025,3)'
.param mc_c_cox_1p0ff='mc_c_cox_1p0ff2*sw_stat_global*cap_mc_skew'
.param mc_c_cox_1p5ff='mc_c_cox_1p5ff2*sw_stat_global*cap_mc_skew'
.param mc_c_cox_2p0ff='mc_c_cox_2p0ff2*sw_stat_global*cap_mc_skew'
.lib 'sm141064.spice' mim_cap
.endl mimcap_statistical
