* Copyright 2022 GlobalFoundries PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.

*******************************************************************************
* Document No.      : SM-BB-000149
* Revision          : 1
* Process Name      : 0.18um MCU 10V high voltage process
* Process ID        : TH18300G1A
*					  TH18300G4A
* Wafer ID          : TNL4435202 (10V LDNMOS & LDPMOS)
************************************************************************************************
* Models included in this release :
*
*      ModelName          Description
*      ---------          -----------
*      nmos_10p0_asym     BSIM4 based HV subcircuit model for 10V LDNMOS (*)
*      pmos_10p0_asym     BSIM4 based HV subcircuit model for 10V LDPMOS (*)
************************************************************************************************

.options parser model_binning=true

.lib typical
.param nmos_10p0_asym_dtox=0
.param nmos_10p0_asym_dxl=0
.param nmos_10p0_asym_dxw=0
.param nmos_10p0_asym_dvth0=0
.param nmos_10p0_asym_drdsw=1
.param nmos_10p0_asym_drdrift=1
.param nmos_10p0_asym_dvsat=1
.param nmos_10p0_asym_du0=1
.param nmos_10p0_asym_dcgs=1
.param nmos_10p0_asym_dcgd=1
.param nmos_10p0_asym_dcjs=1
.param nmos_10p0_asym_dcjd=1
.param pmos_10p0_asym_dtox=0
.param pmos_10p0_asym_dxl=0
.param pmos_10p0_asym_dxw=0
.param pmos_10p0_asym_dvth0=0
.param pmos_10p0_asym_drdsw=1
.param pmos_10p0_asym_drdrift=1
.param pmos_10p0_asym_dvsat=1
.param pmos_10p0_asym_du0=1
.param pmos_10p0_asym_dcgs=1
.param pmos_10p0_asym_dcgd=1
.param pmos_10p0_asym_dcjs=1
.param pmos_10p0_asym_dcjd=1
.lib smbb000149.spice nmos_10p0_asym_t
.lib smbb000149.spice pmos_10p0_asym_t
.lib smbb000149.spice noise_corner
.endl typical

.lib ss
.param nmos_10p0_asym_dtox=8e-10
.param nmos_10p0_asym_dxl=6e-008
.param nmos_10p0_asym_dxw=-3.46e-8
.param nmos_10p0_asym_dvth0=0.112
.param nmos_10p0_asym_drdsw=1.2
.param nmos_10p0_asym_drdrift=1.271
.param nmos_10p0_asym_dvsat=0.926
.param nmos_10p0_asym_du0=0.95
.param nmos_10p0_asym_dcgs=1.1
.param nmos_10p0_asym_dcgd=1.2
.param nmos_10p0_asym_dcjs=1.1
.param nmos_10p0_asym_dcjd=1.2
.param pmos_10p0_asym_dtox=8e-10
.param pmos_10p0_asym_dxl=9.914e-008
.param pmos_10p0_asym_dxw=-1e-7
.param pmos_10p0_asym_dvth0=-0.0936
.param pmos_10p0_asym_drdsw=1.11
.param pmos_10p0_asym_drdrift=1.144
.param pmos_10p0_asym_dvsat=0.91
.param pmos_10p0_asym_du0=0.964
.param pmos_10p0_asym_dcgs=1.1
.param pmos_10p0_asym_dcgd=1.2
.param pmos_10p0_asym_dcjs=1.1
.param pmos_10p0_asym_dcjd=1.2
.lib smbb000149.spice nmos_10p0_asym_t
.lib smbb000149.spice pmos_10p0_asym_t
.lib smbb000149.spice noise_corner
.endl ss

.lib ff
.param nmos_10p0_asym_dtox=-8e-10
.param nmos_10p0_asym_dxl=-6e-008
.param nmos_10p0_asym_dxw=3.46e-8
.param nmos_10p0_asym_dvth0=-0.10388
.param nmos_10p0_asym_drdsw=0.868
.param nmos_10p0_asym_drdrift=0.8245
.param nmos_10p0_asym_dvsat=1.033
.param nmos_10p0_asym_du0=1.04
.param nmos_10p0_asym_dcgs=0.9
.param nmos_10p0_asym_dcgd=0.8
.param nmos_10p0_asym_dcjs=0.9
.param nmos_10p0_asym_dcjd=0.8
.param pmos_10p0_asym_dtox=-8e-10
.param pmos_10p0_asym_dxl=-6.804e-008
.param pmos_10p0_asym_dxw=8.46e-8
.param pmos_10p0_asym_dvth0=0.099
.param pmos_10p0_asym_drdsw=0.91
.param pmos_10p0_asym_drdrift=0.89
.param pmos_10p0_asym_dvsat=1.06
.param pmos_10p0_asym_du0=1.03
.param pmos_10p0_asym_dcgs=0.9
.param pmos_10p0_asym_dcgd=0.8
.param pmos_10p0_asym_dcjs=0.9
.param pmos_10p0_asym_dcjd=0.8
.lib smbb000149.spice nmos_10p0_asym_t
.lib smbb000149.spice pmos_10p0_asym_t
.lib smbb000149.spice noise_corner
.endl ff

.lib sf
.param nmos_10p0_asym_dtox=0
.param nmos_10p0_asym_dxl=5.024e-008
.param nmos_10p0_asym_dxw=0
.param nmos_10p0_asym_dvth0=0.068
.param nmos_10p0_asym_drdsw=1.2
.param nmos_10p0_asym_drdrift=1.156
.param nmos_10p0_asym_dvsat=0.928
.param nmos_10p0_asym_du0=0.97
.param nmos_10p0_asym_dcgs=1.07
.param nmos_10p0_asym_dcgd=1.14
.param nmos_10p0_asym_dcjs=1.07
.param nmos_10p0_asym_dcjd=1.14
.param pmos_10p0_asym_dtox=0
.param pmos_10p0_asym_dxl=-7.004e-008
.param pmos_10p0_asym_dxw=0
.param pmos_10p0_asym_dvth0=0.057672
.param pmos_10p0_asym_drdsw=0.91
.param pmos_10p0_asym_drdrift=0.92
.param pmos_10p0_asym_dvsat=1.012
.param pmos_10p0_asym_du0=1.03
.param pmos_10p0_asym_dcgs=0.93
.param pmos_10p0_asym_dcgd=0.86
.param pmos_10p0_asym_dcjs=0.93
.param pmos_10p0_asym_dcjd=0.86
.lib smbb000149.spice nmos_10p0_asym_t
.lib smbb000149.spice pmos_10p0_asym_t
.lib smbb000149.spice noise_corner
.endl sf

.lib fs
.param nmos_10p0_asym_dtox=0
.param nmos_10p0_asym_dxl=-5.02e-008
.param nmos_10p0_asym_dxw=0
.param nmos_10p0_asym_dvth0=-0.058169
.param nmos_10p0_asym_drdsw=0.868
.param nmos_10p0_asym_drdrift=0.89748
.param nmos_10p0_asym_dvsat=1.045
.param nmos_10p0_asym_du0=1.034
.param nmos_10p0_asym_dcgs=0.93
.param nmos_10p0_asym_dcgd=0.86
.param nmos_10p0_asym_dcjs=0.93
.param nmos_10p0_asym_dcjd=0.86
.param pmos_10p0_asym_dtox=0
.param pmos_10p0_asym_dxl=9.414e-008
.param pmos_10p0_asym_dxw=0
.param pmos_10p0_asym_dvth0=-0.056
.param pmos_10p0_asym_drdsw=1.11
.param pmos_10p0_asym_drdrift=1.06
.param pmos_10p0_asym_dvsat=0.989
.param pmos_10p0_asym_du0=0.97
.param pmos_10p0_asym_dcgs=1.07
.param pmos_10p0_asym_dcgd=1.14
.param pmos_10p0_asym_dcjs=1.07
.param pmos_10p0_asym_dcjd=1.14
.lib smbb000149.spice nmos_10p0_asym_t
.lib smbb000149.spice pmos_10p0_asym_t
.lib smbb000149.spice noise_corner
.endl fs

.lib statistical
.param mc_vsat2_10v='agauss(0,1,3)'
.param mc_rd_10v_2='agauss(0,1,3)'
.param mc_u0_10v_2='agauss(0,1,3)'
.param mc_cgol_10v_2='agauss(0,1,3)'
.param mc_vsatn2_10v='agauss(0,1,3)'
.param mc_rdn_10v_2='agauss(0,1,3)'
.param mc_u0n_10v_2='agauss(0,1,3)'
.param mc_cgoln_10v_2='agauss(0,1,3)'
.param mc_vsatp2_10v='agauss(0,1,3)'
.param mc_u0p2_10v='agauss(0,1,3)'
.param mc_rdp_10v_2='agauss(0,1,3)'
.param mc_cgolp_10v_2='agauss(0,1,3)'
.param mc_vsat_10v='mc_vsat2_10v'
.param mc_rd_10v='mc_rd_10v_2'
.param mc_u0_10v='mc_u0_10v_2'
.param mc_cgol_10v='mc_cgol_10v_2'
.param mc_vsatn_10v='mc_vsatn2_10v'
.param mc_rdn_10v='mc_rdn_10v_2'
.param mc_u0n_10v='mc_u0n_10v_2'
.param mc_cgoln_10v='mc_cgoln_10v_2'
.param mc_vsatp_10v='mc_vsatp2_10v'
.param mc_u0p_10v='mc_u0p2_10v'
.param mc_rdp_10v='mc_rdp_10v_2'
.param mc_cgolp_10v='mc_cgolp_10v_2'
.param nmos_10p0_asym_sig_vth='0.01675*(0.7*mc_sig_vth+0.7*mc_sig_vthn)*sw_stat_global*mc_skew'
.param nmos_10p0_asym_dtox='7.2e-11*(0.77*mc_toxe+0.63*mc_toxen)*sw_stat_global*mc_skew'
.param nmos_10p0_asym_dxl='5.3e-9*(0.71*mc_xl+0.69*mc_xln)*sw_stat_global*mc_skew'
.param nmos_10p0_asym_dxw='3.25e-8*(0.77*mc_xw+0.63*mc_xwn)*sw_stat_global*mc_skew'
.param nmos_10p0_asym_dvth0='nmos_10p0_asym_sig_vth'
.param nmos_10p0_asym_drdsw='(1+0.093*(0.77*mc_rd_10v+0.63*mc_rdn_10v)*sw_stat_global*mc_skew)'
.param nmos_10p0_asym_drdrift='(1+0.037*(0.77*mc_rd_10v+0.63*mc_rdn_10v)*sw_stat_global*mc_skew)'
.param nmos_10p0_asym_dvsat='(1+0.028*(0.77*mc_vsat_10v+0.63*mc_vsatn_10v)*sw_stat_global*mc_skew)'
.param nmos_10p0_asym_du0='(1+0.0157*(0.7*mc_u0_10v+0.7*mc_u0n_10v)*sw_stat_global*mc_skew)'
.param nmos_10p0_asym_dcgs='(1+(12e-3*mc_cgol_10v+12e-3*mc_cgoln_10v)*sw_stat_global*mc_skew)'
.param nmos_10p0_asym_dcgd='(1+(24e-3*mc_cgol_10v+24e-3*mc_cgoln_10v)*sw_stat_global*mc_skew)'
.param nmos_10p0_asym_dcjs='(1+(12e-3*mc_cgol_10v+12e-3*mc_cgoln_10v)*sw_stat_global*mc_skew)'
.param nmos_10p0_asym_dcjd='(1+(24e-3*mc_cgol_10v+24e-3*mc_cgoln_10v)*sw_stat_global*mc_skew)'
.param pmos_10p0_asym_sig_dvth1='0.01692*(-0.7*mc_sig_vth+0.7*mc_sig_vthp)*sw_stat_global*mc_skew'
.param pmos_10p0_asym_dtox='7.143e-11*(0.77*mc_toxe+0.63*mc_toxep)*sw_stat_global*mc_skew'
.param pmos_10p0_asym_dxl='1.7e-8*(0.71*mc_xl+0.69*mc_xlp)*sw_stat_global*mc_skew'
.param pmos_10p0_asym_dxw='7.4e-8*(0.77*mc_xw+0.63*mc_xwp)*sw_stat_global*mc_skew'
.param pmos_10p0_asym_dvth0='pmos_10p0_asym_sig_dvth1'
.param pmos_10p0_asym_drdsw='(1+0.085*(0.77*mc_rd_10v+0.63*mc_rdp_10v)*sw_stat_global*mc_skew)'
.param pmos_10p0_asym_drdrift='(1+0.032*(0.77*mc_rd_10v+0.63*mc_rdp_10v)*sw_stat_global*mc_skew)'
.param pmos_10p0_asym_dvsat='(1+0.032*(0.77*mc_vsat_10v+0.63*mc_vsatp_10v)*sw_stat_global*mc_skew)'
.param pmos_10p0_asym_du0='(1+0.0097*(0.7*mc_u0_10v+0.7*mc_u0p_10v)*sw_stat_global*mc_skew)'
.param pmos_10p0_asym_dcgs='(1+(12e-3*mc_cgol_10v+12e-3*mc_cgolp_10v)*sw_stat_global*mc_skew)'
.param pmos_10p0_asym_dcgd='(1+(24e-3*mc_cgol_10v+24e-3*mc_cgolp_10v)*sw_stat_global*mc_skew)'
.param pmos_10p0_asym_dcjs='(1+(12e-3*mc_cgol_10v+12e-3*mc_cgolp_10v)*sw_stat_global*mc_skew)'
.param pmos_10p0_asym_dcjd='(1+(24e-3*mc_cgol_10v+24e-3*mc_cgolp_10v)*sw_stat_global*mc_skew)'
.lib smbb000149.spice nmos_10p0_asym_t
.lib smbb000149.spice pmos_10p0_asym_t
.lib smbb000149.spice noise_corner
.endl statistical

.lib noise_corner
.param nmos_10p0_asym_noia='(fnoicor==0)*1.1021e42+(fnoicor==1)*2.5852e42'
.param nmos_10p0_asym_noib='(fnoicor==0)*2.8476e24+(fnoicor==1)*6.5096e+024'
.param nmos_10p0_asym_noic='(fnoicor==0)*8.75+(fnoicor==1)*8.75'
.param pmos_10p0_asym_noia='(fnoicor==0)*2.9073e+041+(fnoicor==1)*1.7073e+042'
.param pmos_10p0_asym_noib='(fnoicor==0)*8.0736e+025+(fnoicor==1)*2.4523e+026'
.param pmos_10p0_asym_noic='(fnoicor==0)*12780+(fnoicor==1)*12780'
.endl noise_corner

.lib nmos_10p0_asym_t
.subckt nmos_10p0_asym d g s b params: w=25e-6 l=0.6e-6 ad='w*1.48e-6' pd='2*(1.48e-6+w)' as='w*0.48e-6' ps='(w+0.48e-6)*2' nrd=0 nrs=0 nf=1 dtemp=0 sa=0 sb=0 sd=0 par=1
.param rdrift1=1.5433e3
.param wa=-1.6705e-8
.param rd=0.17322
.param ra=4.631e-3
.param rb=1.1181
.param lb=-1.0648e-6
.param wb=-2.8512e-7
.param trx1=2.8643e-3
.param trx2=1.0098e-5
.param trth1=5.5e-4
.param trth2=0
.param cgdl_d2=5.0343e-10
.param toxep=1.376e-8
.param lcgd_d2=6.4774e-10
.param cgdv_d=1.0253
.param cgd_val=0.20473
.param cgsl_s=1.2929e-10
.param lcgs=2.9695e-8
.param cgs_slope=4.0853
.param cgs_vth=0.10612
.param cgs_factor=0.9
.param vthd=4.18986e-2
.param cgd_vthd=0.31232
.param cgb_slope=1.0158
.param cgb_vth=0.82325
.param cgb_amp=1.3591e-9
.param cgb_min=7.4448e-10
.param cgb_power=2.5552
.param lcgd_d=1.4497e-7
.param polar_d=-1.0276e-3
.param polard_min=7.05
.param polar_s=-0.35192
.param polars_min=4.2
.param cgs_factor2=1
.param cgdv_d2=-2.1473
.param cgdl_d=1.3222e-11
.param cgs_vth1=0.20635
.param cgds_fixed='3.9*8.854e-12/toxep'
rdrift d d2 tc1='trx1' tc2='trx2' m='nf' r='(rdrift1*nmos_10p0_asym_drdrift)*1.2e-6/(w/nf-wa)'
rd2 d2 d1 m='nf' r='max(1e-2,(rd*nmos_10p0_asym_drdsw*(1+trth1*(temp+dtemp-25)+trth2*(temp+dtemp-25)*(temp+dtemp-25)))/(w/nf-wb)*(tanh(ra*(v(d,s)-rb*(l-lb)/(0.6e-6-lb)))))'
m0 d1 g s b nmos_10p0_asym_core ad='ad' as='as' l='l' nf='nf' nrd='nrd' nrs='nrs' pd='pd' ps='ps' sa='sa' sb='sb' sd='sd' w='w'
c1_gd g d c='nmos_10p0_asym_dcgd*(cgds_fixed*w*lcgd_d+exp(polar_d*min(max(v(d,s)-vthd,0),polard_min))*cgdl_d*w*(1+tanh(cgdv_d/(1+cgd_val*max(v(d,g),0))*(v(g,d1)+cgd_vthd*(1+cgdv_d2*v(d,d1))-nmos_10p0_asym_dvth0))))'
c1_gd2 g d1 c='nmos_10p0_asym_dcgd*(cgds_fixed*w*lcgd_d2+cgdl_d2*w*(1+tanh(cgdv_d/(1+cgd_val*max(v(d,g),0))*(v(g,d1)+cgd_vthd*(1+cgdv_d2*v(d,d1))-nmos_10p0_asym_dvth0))))'
c2_gs g s c='nmos_10p0_asym_dcgs*(cgds_fixed*w*lcgs+cgsl_s*w*(1-tanh(cgs_slope*(v(s,g)+cgs_vth)))*(1+cgs_factor/(1+cgs_factor2*exp(-v(g,d1)-cgs_vth1))*(1-exp(polar_s*min(max(v(d1,s)-vthd,0),polars_min)))))'
c3_gb g b c='(cgb_min+cgb_amp/(1+(1/pow(max(1e-3,cgb_slope*(v(b,g)-cgb_vth+nmos_10p0_asym_dvth0)),cgb_power))))*w'
.model nmos_10p0_asym_core.1 nmos a0=1.0212 a1=-0.065307 a2=0.94 acde=0.54775 acnqsmod=0 agidl=5.7877e-16 ags=0.13804 alpha0=-2.5481e-7 alpha1=0.59769 at=3.3e4 b0=6.48e-6 b1=5.9519e-5 beta0=37.485 bgidl=1.171e9 binunit=1 bvd=14.5 bvs=11 capmod=2 cdsc=1.1424e-5 cdscb=2.4894e-6 cdscd=0 cgbo=1e-13 cgdl=0 cgdo=0 cgidl=0.228 cgsl=0 cgso=0 cit=0 cjd='1.4914e-4*nmos_10p0_asym_dcjd' cjs='9.5e-4*nmos_10p0_asym_dcjs' cjswd='5.8719e-10*nmos_10p0_asym_dcjd' cjswgd='5.8719e-10*nmos_10p0_asym_dcjd' cjswgs='1.33e-10*nmos_10p0_asym_dcjs' cjsws='1.33e-10*nmos_10p0_asym_dcjs' ckappad=0.6 ckappas=0.6 delta=0.01 diomod=2 dlc=1.723e-7 drout=0.45 dsub=0.56 dvt0=0.09762 dvt0w=3.4488 dvt1=0.021131 dvt1w=9.5865e4 dvt2=-0.046683 dvt2w=0.034426 dvtp0=0 dvtp1=0 dwb=-3.3647e-8 dwg=-2.9807e-8 ef=1.0914 egidl=0.0968 em=4.1e7 epsrox=3.9 eta0=0.039833 etab=-1.2928 fnoimod=1 geomod=0 igbmod=0 igcmod=0 jsd=1.6119e-6 jss=6.88e-7 jswd=4.824e-12 jswgd=4.824e-12 jswgs=4.88e-13 jsws=4.88e-13 jtsd=1.4513e-4 k1=0.9621 k2=-7.2357e-3 k3=13.237 k3b=0.25485 keta=-0.01362 kt1=-0.42425 kt1l=-1.8892e-8 kt2=-0.060553 la0=-0.55504 lags=0 lat=0 lbeta0=-11.164 lint=0 lk1=0 lk2=0 lketa=-3.3807e-3 ll=0 lln=1 lmax=20.01e-6 lmin=6e-7 lnfactor=6.48e-7 lnoff=1 lpe0=1.0439e-6 lpeb=6.2517e-7 lu0='5.2003e-3*nmos_10p0_asym_du0' lua=4.2194e-10 lua1=0 lub=-1.9302e-18 lub1=0 luc=-4.7702e-11 lute=0.045577 lvsat='9844*nmos_10p0_asym_dvsat' lvth0=0 lw=0 lwl=0 lwn=1 minv=0 mjd=0.30525 mjs=0.296 mjswd=0.21757 mjswgd=0.21757 mjswgs=0.01 mjsws=0.01 mobmod=0 moin=16.92 ndep=1.7e17 nfactor=0.90694 ngate=2.9861e21 njd=1 njs=1.0541 noff=1.9257 noia='nmos_10p0_asym_noia' noib='nmos_10p0_asym_noib' noic='nmos_10p0_asym_noic' nsd=1e20 paramchk=1 pat=-9e3 pbd=0.43905 pbeta0=-0.645 pbs=0.606 pbswd=0.48991 pbswgd=0.48991 pbswgs=0.48 pbsws=0.48 pclm=0.02794 pdiblc1=0.46226 pdiblc2=1.092e-4 pdiblcb=-5e-3 permod=1 phin=0 pkt1=0 pkt2=-0.09625 pprt=0 pprwb=0 pprwg=0 prdsw=0 prt=200 prwb=0.81 prwg=0.037838 pscbe1=4.9654e8 pscbe2=1.6381e-7 pu0='3.9064e-3*nmos_10p0_asym_du0' pua=0 pua1=0 pub=-6.8e-19 pub1=0 puc=-6.8588e-11 pute=0.17695 pvag=0.9 pvsat=-3.168e3 pvth0=0.19879 rbodymod=0 rdsmod=0 rdsw='200*nmos_10p0_asym_drdsw' rdswmin=500 rsh=7 tcj=1.65e-3 tcjsw=1.61e-3 tcjswg=1.61e-3 tempmod=0 tnoimod=0 tnom=25 toxe='1.398e-8+nmos_10p0_asym_dtox' tpb=2.11e-3 tpbsw=1.9e-3 tpbswg=1.9e-3 trnqsmod=0 u0='0.0486*nmos_10p0_asym_du0' ua=-1.05e-10 ua1=3.2446e-9 ub=3.0678e-18 ub1=-4.2148e-18 uc=1.0312e-10 uc1=-7.2993e-11 ute=-1.3028 vfb=-0.55 voff=-0.092552 voffcv=-0.038 voffl=-1.4059e-8 vsat='7.9784e4*nmos_10p0_asym_dvsat' vth0='0.653+nmos_10p0_asym_dvth0' vtsd=2.16 w0=1e-6 wags=-0.012 wbeta0=2.034 wint=0 wk3=0 wkt1=0 wl=0 wln=1 wmax=50.01e-6 wmin=4e-6 wr=1 wu0='-0.020672*nmos_10p0_asym_du0' wvsat=0 wvth0=0 ww=0 wwl=0 wwn=1 xj=1.5e-7 xjbvd=1 xjbvs=1 xl='0+nmos_10p0_asym_dxl' xpart=1 xtid=3 xtis=3 xtsd=0.63818 xw='0+nmos_10p0_asym_dxw' level=14
.ends nmos_10p0_asym
.endl nmos_10p0_asym_t

.lib pmos_10p0_asym_t
.subckt pmos_10p0_asym d g s b params: w=2.5e-5 l=6e-7 dtemp=0 nf=1 ad='(w*1.78e-6)' pd='2*(w+1.78e-6)' as='w*0.48e-6' ps='(w+0.48e-6)*2' nrd=0 nrs=0 sa=0 sb=0 sd=0 par=1
.param rdrift=5.751e-3
.param rd=0.94645
.param ra=1.1954e-3
.param rb=1.5957
.param lb=6.78e-6
.param wa=-6.5504e-7
.param wb=4.1955e-8
.param trx1=2.836e-3
.param trx2=7.4236e-6
.param trd1=-3.7522e-3
.param cgdl_d2=4.3795e-10
.param toxep=1.568e-8
.param lcgd_d2=6.4774e-10
.param cgdv_d=1.0253
.param cgd_val=0.20473
.param cgsl_s=1.2929e-11
.param lcgs=6.4247e-9
.param cgs_slope=0.81706
.param cgs_vth=0.021224
.param cgs_factor=0.9
.param vthd=4.18986e-2
.param cgd_vthd=0.31232
.param cgb_slope=1.0219
.param cgb_vth=0.89948
.param cgb_amp=9.9049e-10
.param cgb_min=3.2564e-11
.param cgb_power=2.5552
.param lcgd_d=1.4497e-7
.param polar_d=-4.1926e-4
.param polard_min=7.05
.param polar_s=-0.35192
.param polars_min=4.2
.param cgs_factor2=1
.param cgdv_d2=-1.2197
.param cgdl_d=1.6046e-11
.param cgs_vth1=0.13041
.param cgds_fixed='3.9*8.854e-12/toxep'
rd1 d d2 tc1='trx1' tc2='trx2' m='nf' r='(rdrift*pmos_10p0_asym_drdrift)/(w/nf-wa)'
rd2 d2 d1 m='nf' r='max(0.1,(rd*pmos_10p0_asym_drdsw*(1+trd1*(temp+dtemp-25))/(w/nf-wb)*(tanh(ra*(v(s,d)-rb*(l-lb)/(0.6e-6-lb))))))'
m0 d1 g s b pmos_10p0_asym_core ad='ad' as='as' l='l' nf='nf' nrd='nrd' nrs='nrs' pd='pd' ps='ps' sa='sa' sb='sb' sd='sd' w='w'
c1_gd g d c='pmos_10p0_asym_dcgd*(cgds_fixed*w*lcgd_d+exp(polar_d*min(max(-v(d,s)-vthd,0),polard_min))*cgdl_d*w*(1+tanh(cgdv_d/(1+cgd_val*max(-v(d,g),0))*(-v(g,d1)+cgd_vthd*(1+cgdv_d2*-v(d,d1))-pmos_10p0_asym_dvth0))))'
c1_gd2 g d1 c='pmos_10p0_asym_dcgd*(cgds_fixed*w*lcgd_d2+cgdl_d2*w*(1+tanh(cgdv_d/(1+cgd_val*max(-v(d,g),0))*(-v(g,d1)+cgd_vthd*(1+cgdv_d2*-v(d,d1))-pmos_10p0_asym_dvth0))))'
c2_gs g s c='pmos_10p0_asym_dcgs*(cgds_fixed*w*lcgs+cgsl_s*w*(1-tanh(cgs_slope*(-v(s,g)+cgs_vth)))*(1+cgs_factor/(1+cgs_factor2*exp(v(g,d1)-cgs_vth1))*(1-exp(polar_s*min(max(-v(d1,s)-vthd,0),polars_min)))))'
c3_gb g b c='(cgb_min+cgb_amp/(1+(1/pow(max(1e-3,cgb_slope*(-v(b,g)-cgb_vth+pmos_10p0_asym_dvth0)),cgb_power))))*w'
.model pmos_10p0_asym_core.1 pmos a0=1.1348 a1=-0.07052 a2=1 acde=1 acnqsmod=0 agidl=3.7498e-17 ags=0.0834 aigbacc=0.43 aigbinv=0.35 aigc=0.43 aigsd=0.43 alpha0=7.0634e-8 alpha1=0.14712 at=3.96e3 b0=0 b1=0 beta0=66.68 bgidl=1.196e8 bigbacc=0.054 bigbinv=0.03 bigc=0.054 bigsd=0.054 binunit=2 bvd=14.5 bvs=10.5 capmod=2 cdsc=4.248e-4 cdscb=6e-5 cdscd=0 cgbo=0 cgdl=0 cgdo=0 cgidl=0.5 cgsl=0 cgso=0 cigbacc=0.075 cigbinv=6e-3 cigc=0.075 cigsd=0.075 cit=0 cjd='3.2124e-4*pmos_10p0_asym_dcjd' cjs='9.12e-4*pmos_10p0_asym_dcjs' cjswd='5.4659e-10*pmos_10p0_asym_dcjd' cjswgd='5.4659e-10*pmos_10p0_asym_dcjd' cjswgs='1.4649e-10*pmos_10p0_asym_dcjs' cjsws='1.4649e-10*pmos_10p0_asym_dcjs' ckappad=0.6 ckappas=0.6 clc=1e-7 cle=0.6 delta=0.01 diomod=0 dlc=5.0579e-8 drout=0.56 dsub=0.56 dvt0=4.0503 dvt0w=0 dvt1=0.16044 dvt1w=2.7518e4 dvt2=-0.038473 dvt2w=-0.032 dvtp0=0 dvtp1=0 dwb=0 dwg=1.0544e-8 ef=1.1237 egidl=0.8 eigbinv=1.1 em=4.1e7 epsrox=3.9 eta0=0.08 etab=-0.57865 eu=1.67 fnoimod=1 fprout=0 geomod=0 igbmod=0 igcmod=0 jsd=5.2139e-7 jss=2.0867e-7 jswd=1.5e-13 jswgd=1.5e-13 jswgs=1.6088e-13 jsws=1.6088e-13 jtsd=1.0891e-6 k1=1.09 k2=-0.014623 k3=5.4746 k3b=3.8727 keta=-1.504e-3 kt1=-0.45028 kt1l=-4.1552e-8 kt2=-0.05137 la0=-3.8459e-7 lags=0 lbeta0=-2.1875e-6 lint=0 lketa=-2.0415e-8 ll=0 llpe0=0 lmax=20.01e-6 lmin=6e-7 lnoff=1.2657e-6 lpe0=2.814e-7 lpeb=3.068e-7 lu0='2.7385e-9*pmos_10p0_asym_du0' lua=1.2893e-16 lua1=0 lub=0 lub1=-2.0019e-25 luc=5.88e-17 luc1=0 lute=-1.1751e-7 lwl=0 minv=0 mjd=0.31113 mjs=0.32713 mjswd=0.39816 mjswgd=0.39816 mjswgs=0.056777 mjsws=0.056777 mobmod=0 moin=11.1 ndep=1.7e17 nfactor=1.096 ngate=1e20 nigbacc=1 nigbinv=3 nigc=1 noff=1.8144 noia='pmos_10p0_asym_noia' noib='pmos_10p0_asym_noib' noic='pmos_10p0_asym_noic' nsd=1e20 ntox=1 pags=6.4229e-13 paramchk=1 pbd=0.63391 pbeta0=0 pbs=0.76836 pbswd=0.77752 pbswgd=0.77752 pbswgs=0.5 pbsws=0.5 pclm=0.37315 pdiblc1=0.09466 pdiblc2=5.586e-8 pdiblcb=0 pdits=0 pditsd=0 pditsl=0 pdvt0=-2.3525e-12 pdvt1=0 permod=1 phin=0.061992 pigcd=1 pk2=-9.04e-14 pketa=-7.5094e-014 pkt1=0 pkt2=-1.1e-13 plpe0=0 poxedge=1 prt=0 prwb=1.24 prwg=1 pscbe1=5.9843e8 pscbe2=9.3757e-8 pu0='-2e-15*pmos_10p0_asym_du0' pua=6.315e-22 pute=1.0911e-13 pvag=1.2 pvsat=0 pvth0=1.44e-14 rbodymod=0 rdsmod=0 rdsw='200*pmos_10p0_asym_drdsw' rdswmin=0 rdw=100 rdwmin=0 rsh=5.6 rshg=0.4 rsw=100 rswmin=0 tempmod=0 tnoimod=0 toxe='1.568e-8+pmos_10p0_asym_dtox' trnqsmod=0 u0='0.013723*pmos_10p0_asym_du0' ua=1.26e-9 ua1=5e-10 ub=7.2608e-19 ub1=-2.2324e-18 uc=-4.5217e-11 uc1=-3.0912e-11 ute=-1.245 vbm=-3 vfb=-1 vfbcv=-1 voff=-0.08768 voffcv=-3.8635e-3 voffl=0 vsat='71505*pmos_10p0_asym_dvsat' vth0='-0.888+pmos_10p0_asym_dvth0' vtsd=2.44 w0=3.24e-6 wags=6.5664e-9 wbeta0=4.86e-6 wdvt0=0 wdvt1=0 wint=0 wk2=0 wketa=2.68e-008 wkt1=0 wlpe0=-3.5894e-13 wmax=50.01e-6 wmin=4e-6 wr=1 wu0='-7e-10*pmos_10p0_asym_du0' wute=-4e-8 wvsat=0 wvth0=0 ww=0 wwl=0 xj=1.5e-7 xjbvd=1 xjbvs=1 xl='0+pmos_10p0_asym_dxl' xtsd=0.92538 xw='0+pmos_10p0_asym_dxw' level=14
.ends pmos_10p0_asym
.endl pmos_10p0_asym_t
